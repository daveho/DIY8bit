// 800x600 SVGA timing constants

localparam H_VISIBLE_END     = 16'd799;
localparam H_FRONT_PORCH_END = 16'd839;
localparam H_SYNC_PULSE_END  = 16'd967;
localparam H_BACK_PORCH_END  = 16'd1055;

localparam V_VISIBLE_END     = 16'd599;
localparam V_FRONT_PORCH_END = 16'd600;
localparam V_SYNC_PULSE_END  = 16'd604;
localparam V_BACK_PORCH_END  = 16'd627;

// vim:ft=verilog:
