vramDataLower[12'd0] = 8'd31;
vramDataLower[12'd1] = 8'd199;
vramDataLower[12'd2] = 8'd202;
vramDataLower[12'd3] = 8'd87;
vramDataLower[12'd4] = 8'd252;
vramDataLower[12'd5] = 8'd87;
vramDataLower[12'd6] = 8'd200;
vramDataLower[12'd7] = 8'd151;
vramDataLower[12'd8] = 8'd220;
vramDataLower[12'd9] = 8'd121;
vramDataLower[12'd10] = 8'd220;
vramDataLower[12'd11] = 8'd121;
vramDataLower[12'd12] = 8'd183;
vramDataLower[12'd13] = 8'd121;
vramDataLower[12'd14] = 8'd214;
vramDataLower[12'd15] = 8'd121;
vramDataLower[12'd16] = 8'd223;
vramDataLower[12'd17] = 8'd151;
vramDataLower[12'd18] = 8'd223;
vramDataLower[12'd19] = 8'd151;
vramDataLower[12'd20] = 8'd188;
vramDataLower[12'd21] = 8'd151;
vramDataLower[12'd22] = 8'd214;
vramDataLower[12'd23] = 8'd247;
vramDataLower[12'd24] = 8'd202;
vramDataLower[12'd25] = 8'd247;
vramDataLower[12'd26] = 8'd210;
vramDataLower[12'd27] = 8'd151;
vramDataLower[12'd28] = 8'd202;
vramDataLower[12'd29] = 8'd247;
vramDataLower[12'd30] = 8'd210;
vramDataLower[12'd31] = 8'd247;
vramDataLower[12'd32] = 8'd200;
vramDataLower[12'd33] = 8'd135;
vramDataLower[12'd34] = 8'd164;
vramDataLower[12'd35] = 8'd120;
vramDataLower[12'd36] = 8'd210;
vramDataLower[12'd37] = 8'd135;
vramDataLower[12'd38] = 8'd210;
vramDataLower[12'd39] = 8'd135;
vramDataLower[12'd40] = 8'd210;
vramDataLower[12'd41] = 8'd135;
vramDataLower[12'd42] = 8'd16;
vramDataLower[12'd43] = 8'd135;
vramDataLower[12'd44] = 8'd16;
vramDataLower[12'd45] = 8'd120;
vramDataLower[12'd46] = 8'd230;
vramDataLower[12'd47] = 8'd135;
vramDataLower[12'd48] = 8'd30;
vramDataLower[12'd49] = 8'd135;
vramDataLower[12'd50] = 8'd209;
vramDataLower[12'd51] = 8'd135;
vramDataLower[12'd52] = 8'd16;
vramDataLower[12'd53] = 8'd120;
vramDataLower[12'd54] = 8'd210;
vramDataLower[12'd55] = 8'd120;
vramDataLower[12'd56] = 8'd228;
vramDataLower[12'd57] = 8'd120;
vramDataLower[12'd58] = 8'd30;
vramDataLower[12'd59] = 8'd120;
vramDataLower[12'd60] = 8'd210;
vramDataLower[12'd61] = 8'd120;
vramDataLower[12'd62] = 8'd16;
vramDataLower[12'd63] = 8'd135;
vramDataLower[12'd64] = 8'd16;
vramDataLower[12'd65] = 8'd135;
vramDataLower[12'd66] = 8'd16;
vramDataLower[12'd67] = 8'd247;
vramDataLower[12'd68] = 8'd135;
vramDataLower[12'd69] = 8'd120;
vramDataLower[12'd70] = 8'd248;
vramDataLower[12'd71] = 8'd136;
vramDataLower[12'd72] = 8'd0;
vramDataLower[12'd73] = 8'd88;
vramDataLower[12'd74] = 8'd231;
vramDataLower[12'd75] = 8'd136;
vramDataLower[12'd76] = 8'd0;
vramDataLower[12'd77] = 8'd104;
vramDataLower[12'd78] = 8'd17;
vramDataLower[12'd79] = 8'd136;
vramDataLower[12'd80] = 8'd94;
vramDataLower[12'd81] = 8'd200;
vramDataLower[12'd82] = 8'd94;
vramDataLower[12'd83] = 8'd120;
vramDataLower[12'd84] = 8'd252;
vramDataLower[12'd85] = 8'd120;
vramDataLower[12'd86] = 8'd252;
vramDataLower[12'd87] = 8'd120;
vramDataLower[12'd88] = 8'd252;
vramDataLower[12'd89] = 8'd120;
vramDataLower[12'd90] = 8'd252;
vramDataLower[12'd91] = 8'd120;
vramDataLower[12'd92] = 8'd202;
vramDataLower[12'd93] = 8'd120;
vramDataLower[12'd94] = 8'd202;
vramDataLower[12'd95] = 8'd120;
vramDataLower[12'd96] = 8'd202;
vramDataLower[12'd97] = 8'd120;
vramDataLower[12'd98] = 8'd202;
vramDataLower[12'd99] = 8'd120;
vramDataLower[12'd100] = 8'd202;
vramDataLower[12'd101] = 8'd120;
vramDataLower[12'd102] = 8'd31;
vramDataLower[12'd103] = 8'd120;
vramDataLower[12'd104] = 8'd31;
vramDataLower[12'd105] = 8'd120;
vramDataLower[12'd106] = 8'd31;
vramDataLower[12'd107] = 8'd120;
vramDataLower[12'd108] = 8'd31;
vramDataLower[12'd109] = 8'd120;
vramDataLower[12'd110] = 8'd30;
vramDataLower[12'd111] = 8'd120;
vramDataLower[12'd112] = 8'd16;
vramDataLower[12'd113] = 8'd120;
vramDataLower[12'd114] = 8'd16;
vramDataLower[12'd115] = 8'd168;
vramDataLower[12'd116] = 8'd30;
vramDataLower[12'd117] = 8'd168;
vramDataLower[12'd118] = 8'd30;
vramDataLower[12'd119] = 8'd200;
vramDataLower[12'd120] = 8'd214;
vramDataLower[12'd121] = 8'd120;
vramDataLower[12'd122] = 8'd30;
vramDataLower[12'd123] = 8'd120;
vramDataLower[12'd124] = 8'd248;
vramDataLower[12'd125] = 8'd120;
vramDataLower[12'd126] = 8'd193;
vramDataLower[12'd127] = 8'd136;
vramDataLower[12'd128] = 8'd95;
vramDataLower[12'd129] = 8'd152;
vramDataLower[12'd130] = 8'd213;
vramDataLower[12'd131] = 8'd120;
vramDataLower[12'd132] = 8'd197;
vramDataLower[12'd133] = 8'd120;
vramDataLower[12'd134] = 8'd210;
vramDataLower[12'd135] = 8'd120;
vramDataLower[12'd136] = 8'd198;
vramDataLower[12'd137] = 8'd120;
vramDataLower[12'd138] = 8'd164;
vramDataLower[12'd139] = 8'd135;
vramDataLower[12'd140] = 8'd30;
vramDataLower[12'd141] = 8'd135;
vramDataLower[12'd142] = 8'd80;
vramDataLower[12'd143] = 8'd135;
vramDataLower[12'd144] = 8'd150;
vramDataLower[12'd145] = 8'd87;
vramDataLower[12'd146] = 8'd16;
vramDataLower[12'd147] = 8'd135;
vramDataLower[12'd148] = 8'd16;
vramDataLower[12'd149] = 8'd87;
vramDataLower[12'd150] = 8'd126;
vramDataLower[12'd151] = 8'd119;
vramDataLower[12'd152] = 8'd219;
vramDataLower[12'd153] = 8'd126;
vramDataLower[12'd154] = 8'd198;
vramDataLower[12'd155] = 8'd55;
vramDataLower[12'd156] = 8'd16;
vramDataLower[12'd157] = 8'd120;
vramDataLower[12'd158] = 8'd213;
vramDataLower[12'd159] = 8'd120;
vramDataLower[12'd160] = 8'd31;
vramDataLower[12'd161] = 8'd247;
vramDataLower[12'd162] = 8'd31;
vramDataLower[12'd163] = 8'd247;
vramDataLower[12'd164] = 8'd36;
vramDataLower[12'd165] = 8'd119;
vramDataLower[12'd166] = 8'd31;
vramDataLower[12'd167] = 8'd87;
vramDataLower[12'd168] = 8'd24;
vramDataLower[12'd169] = 8'd119;
vramDataLower[12'd170] = 8'd196;
vramDataLower[12'd171] = 8'd247;
vramDataLower[12'd172] = 8'd200;
vramDataLower[12'd173] = 8'd247;
vramDataLower[12'd174] = 8'd202;
vramDataLower[12'd175] = 8'd247;
vramDataLower[12'd176] = 8'd202;
vramDataLower[12'd177] = 8'd247;
vramDataLower[12'd178] = 8'd202;
vramDataLower[12'd179] = 8'd247;
vramDataLower[12'd180] = 8'd202;
vramDataLower[12'd181] = 8'd247;
vramDataLower[12'd182] = 8'd70;
vramDataLower[12'd183] = 8'd247;
vramDataLower[12'd184] = 8'd202;
vramDataLower[12'd185] = 8'd151;
vramDataLower[12'd186] = 8'd212;
vramDataLower[12'd187] = 8'd247;
vramDataLower[12'd188] = 8'd202;
vramDataLower[12'd189] = 8'd247;
vramDataLower[12'd190] = 8'd202;
vramDataLower[12'd191] = 8'd247;
vramDataLower[12'd192] = 8'd16;
vramDataLower[12'd193] = 8'd247;
vramDataLower[12'd194] = 8'd200;
vramDataLower[12'd195] = 8'd87;
vramDataLower[12'd196] = 8'd200;
vramDataLower[12'd197] = 8'd135;
vramDataLower[12'd198] = 8'd202;
vramDataLower[12'd199] = 8'd135;
vramDataLower[12'd200] = 8'd210;
vramDataLower[12'd201] = 8'd152;
vramDataLower[12'd202] = 8'd80;
vramDataLower[12'd203] = 8'd135;
vramDataLower[12'd204] = 8'd202;
vramDataLower[12'd205] = 8'd135;
vramDataLower[12'd206] = 8'd164;
vramDataLower[12'd207] = 8'd120;
vramDataLower[12'd208] = 8'd202;
vramDataLower[12'd209] = 8'd120;
vramDataLower[12'd210] = 8'd181;
vramDataLower[12'd211] = 8'd120;
vramDataLower[12'd212] = 8'd210;
vramDataLower[12'd213] = 8'd120;
vramDataLower[12'd214] = 8'd135;
vramDataLower[12'd215] = 8'd120;
vramDataLower[12'd216] = 8'd145;
vramDataLower[12'd217] = 8'd120;
vramDataLower[12'd218] = 8'd210;
vramDataLower[12'd219] = 8'd120;
vramDataLower[12'd220] = 8'd16;
vramDataLower[12'd221] = 8'd135;
vramDataLower[12'd222] = 8'd85;
vramDataLower[12'd223] = 8'd135;
vramDataLower[12'd224] = 8'd67;
vramDataLower[12'd225] = 8'd87;
vramDataLower[12'd226] = 8'd172;
vramDataLower[12'd227] = 8'd135;
vramDataLower[12'd228] = 8'd31;
vramDataLower[12'd229] = 8'd247;
vramDataLower[12'd230] = 8'd200;
vramDataLower[12'd231] = 8'd135;
vramDataLower[12'd232] = 8'd95;
vramDataLower[12'd233] = 8'd120;
vramDataLower[12'd234] = 8'd214;
vramDataLower[12'd235] = 8'd120;
vramDataLower[12'd236] = 8'd95;
vramDataLower[12'd237] = 8'd120;
vramDataLower[12'd238] = 8'd95;
vramDataLower[12'd239] = 8'd120;
vramDataLower[12'd240] = 8'd95;
vramDataLower[12'd241] = 8'd152;
vramDataLower[12'd242] = 8'd240;
vramDataLower[12'd243] = 8'd136;
vramDataLower[12'd244] = 8'd160;
vramDataLower[12'd245] = 8'd136;
vramDataLower[12'd246] = 8'd175;
vramDataLower[12'd247] = 8'd136;
vramDataLower[12'd248] = 8'd171;
vramDataLower[12'd249] = 8'd136;
vramDataLower[12'd250] = 8'd219;
vramDataLower[12'd251] = 8'd131;
vramDataLower[12'd252] = 8'd255;
vramDataLower[12'd253] = 8'd200;
vramDataLower[12'd254] = 8'd32;
vramDataLower[12'd255] = 8'd72;
vramDataLower[12'd256] = 8'd81;
vramDataLower[12'd257] = 8'd136;
vramDataLower[12'd258] = 8'd149;
vramDataLower[12'd259] = 8'd136;
vramDataLower[12'd260] = 8'd240;
vramDataLower[12'd261] = 8'd136;
vramDataLower[12'd262] = 8'd44;
vramDataLower[12'd263] = 8'd120;
vramDataLower[12'd264] = 8'd140;
vramDataLower[12'd265] = 8'd136;
vramDataLower[12'd266] = 8'd219;
vramDataLower[12'd267] = 8'd128;
vramDataLower[12'd268] = 8'd126;
vramDataLower[12'd269] = 8'd136;
vramDataLower[12'd270] = 8'd0;
vramDataLower[12'd271] = 8'd8;
vramDataLower[12'd272] = 8'd255;
vramDataLower[12'd273] = 8'd232;
vramDataLower[12'd274] = 8'd32;
vramDataLower[12'd275] = 8'd200;
vramDataLower[12'd276] = 8'd214;
vramDataLower[12'd277] = 8'd120;
vramDataLower[12'd278] = 8'd210;
vramDataLower[12'd279] = 8'd120;
vramDataLower[12'd280] = 8'd70;
vramDataLower[12'd281] = 8'd120;
vramDataLower[12'd282] = 8'd253;
vramDataLower[12'd283] = 8'd152;
vramDataLower[12'd284] = 8'd96;
vramDataLower[12'd285] = 8'd152;
vramDataLower[12'd286] = 8'd195;
vramDataLower[12'd287] = 8'd152;
vramDataLower[12'd288] = 8'd30;
vramDataLower[12'd289] = 8'd120;
vramDataLower[12'd290] = 8'd16;
vramDataLower[12'd291] = 8'd120;
vramDataLower[12'd292] = 8'd30;
vramDataLower[12'd293] = 8'd120;
vramDataLower[12'd294] = 8'd17;
vramDataLower[12'd295] = 8'd120;
vramDataLower[12'd296] = 8'd210;
vramDataLower[12'd297] = 8'd120;
vramDataLower[12'd298] = 8'd166;
vramDataLower[12'd299] = 8'd135;
vramDataLower[12'd300] = 8'd253;
vramDataLower[12'd301] = 8'd103;
vramDataLower[12'd302] = 8'd39;
vramDataLower[12'd303] = 8'd135;
vramDataLower[12'd304] = 8'd95;
vramDataLower[12'd305] = 8'd247;
vramDataLower[12'd306] = 8'd126;
vramDataLower[12'd307] = 8'd87;
vramDataLower[12'd308] = 8'd248;
vramDataLower[12'd309] = 8'd55;
vramDataLower[12'd310] = 8'd35;
vramDataLower[12'd311] = 8'd119;
vramDataLower[12'd312] = 8'd67;
vramDataLower[12'd313] = 8'd119;
vramDataLower[12'd314] = 8'd198;
vramDataLower[12'd315] = 8'd55;
vramDataLower[12'd316] = 8'd80;
vramDataLower[12'd317] = 8'd120;
vramDataLower[12'd318] = 8'd16;
vramDataLower[12'd319] = 8'd135;
vramDataLower[12'd320] = 8'd210;
vramDataLower[12'd321] = 8'd183;
vramDataLower[12'd322] = 8'd210;
vramDataLower[12'd323] = 8'd183;
vramDataLower[12'd324] = 8'd210;
vramDataLower[12'd325] = 8'd183;
vramDataLower[12'd326] = 8'd210;
vramDataLower[12'd327] = 8'd183;
vramDataLower[12'd328] = 8'd210;
vramDataLower[12'd329] = 8'd183;
vramDataLower[12'd330] = 8'd210;
vramDataLower[12'd331] = 8'd183;
vramDataLower[12'd332] = 8'd16;
vramDataLower[12'd333] = 8'd151;
vramDataLower[12'd334] = 8'd16;
vramDataLower[12'd335] = 8'd55;
vramDataLower[12'd336] = 8'd202;
vramDataLower[12'd337] = 8'd103;
vramDataLower[12'd338] = 8'd202;
vramDataLower[12'd339] = 8'd103;
vramDataLower[12'd340] = 8'd202;
vramDataLower[12'd341] = 8'd103;
vramDataLower[12'd342] = 8'd202;
vramDataLower[12'd343] = 8'd103;
vramDataLower[12'd344] = 8'd202;
vramDataLower[12'd345] = 8'd231;
vramDataLower[12'd346] = 8'd202;
vramDataLower[12'd347] = 8'd231;
vramDataLower[12'd348] = 8'd80;
vramDataLower[12'd349] = 8'd231;
vramDataLower[12'd350] = 8'd214;
vramDataLower[12'd351] = 8'd183;
vramDataLower[12'd352] = 8'd202;
vramDataLower[12'd353] = 8'd151;
vramDataLower[12'd354] = 8'd209;
vramDataLower[12'd355] = 8'd151;
vramDataLower[12'd356] = 8'd210;
vramDataLower[12'd357] = 8'd183;
vramDataLower[12'd358] = 8'd16;
vramDataLower[12'd359] = 8'd183;
vramDataLower[12'd360] = 8'd202;
vramDataLower[12'd361] = 8'd183;
vramDataLower[12'd362] = 8'd202;
vramDataLower[12'd363] = 8'd55;
vramDataLower[12'd364] = 8'd200;
vramDataLower[12'd365] = 8'd135;
vramDataLower[12'd366] = 8'd209;
vramDataLower[12'd367] = 8'd120;
vramDataLower[12'd368] = 8'd202;
vramDataLower[12'd369] = 8'd135;
vramDataLower[12'd370] = 8'd202;
vramDataLower[12'd371] = 8'd135;
vramDataLower[12'd372] = 8'd16;
vramDataLower[12'd373] = 8'd135;
vramDataLower[12'd374] = 8'd202;
vramDataLower[12'd375] = 8'd135;
vramDataLower[12'd376] = 8'd188;
vramDataLower[12'd377] = 8'd135;
vramDataLower[12'd378] = 8'd248;
vramDataLower[12'd379] = 8'd135;
vramDataLower[12'd380] = 8'd248;
vramDataLower[12'd381] = 8'd135;
vramDataLower[12'd382] = 8'd0;
vramDataLower[12'd383] = 8'd151;
vramDataLower[12'd384] = 8'd235;
vramDataLower[12'd385] = 8'd119;
vramDataLower[12'd386] = 8'd176;
vramDataLower[12'd387] = 8'd119;
vramDataLower[12'd388] = 8'd44;
vramDataLower[12'd389] = 8'd247;
vramDataLower[12'd390] = 8'd200;
vramDataLower[12'd391] = 8'd247;
vramDataLower[12'd392] = 8'd16;
vramDataLower[12'd393] = 8'd247;
vramDataLower[12'd394] = 8'd94;
vramDataLower[12'd395] = 8'd55;
vramDataLower[12'd396] = 8'd210;
vramDataLower[12'd397] = 8'd247;
vramDataLower[12'd398] = 8'd16;
vramDataLower[12'd399] = 8'd247;
vramDataLower[12'd400] = 8'd94;
vramDataLower[12'd401] = 8'd135;
vramDataLower[12'd402] = 8'd94;
vramDataLower[12'd403] = 8'd135;
vramDataLower[12'd404] = 8'd223;
vramDataLower[12'd405] = 8'd135;
vramDataLower[12'd406] = 8'd16;
vramDataLower[12'd407] = 8'd120;
vramDataLower[12'd408] = 8'd95;
vramDataLower[12'd409] = 8'd120;
vramDataLower[12'd410] = 8'd95;
vramDataLower[12'd411] = 8'd152;
vramDataLower[12'd412] = 8'd95;
vramDataLower[12'd413] = 8'd152;
vramDataLower[12'd414] = 8'd218;
vramDataLower[12'd415] = 8'd120;
vramDataLower[12'd416] = 8'd223;
vramDataLower[12'd417] = 8'd135;
vramDataLower[12'd418] = 8'd95;
vramDataLower[12'd419] = 8'd120;
vramDataLower[12'd420] = 8'd230;
vramDataLower[12'd421] = 8'd120;
vramDataLower[12'd422] = 8'd6;
vramDataLower[12'd423] = 8'd136;
vramDataLower[12'd424] = 8'd219;
vramDataLower[12'd425] = 8'd129;
vramDataLower[12'd426] = 8'd182;
vramDataLower[12'd427] = 8'd136;
vramDataLower[12'd428] = 8'd183;
vramDataLower[12'd429] = 8'd152;
vramDataLower[12'd430] = 8'd218;
vramDataLower[12'd431] = 8'd120;
vramDataLower[12'd432] = 8'd210;
vramDataLower[12'd433] = 8'd120;
vramDataLower[12'd434] = 8'd30;
vramDataLower[12'd435] = 8'd120;
vramDataLower[12'd436] = 8'd223;
vramDataLower[12'd437] = 8'd120;
vramDataLower[12'd438] = 8'd248;
vramDataLower[12'd439] = 8'd120;
vramDataLower[12'd440] = 8'd165;
vramDataLower[12'd441] = 8'd136;
vramDataLower[12'd442] = 8'd244;
vramDataLower[12'd443] = 8'd136;
vramDataLower[12'd444] = 8'd214;
vramDataLower[12'd445] = 8'd152;
vramDataLower[12'd446] = 8'd30;
vramDataLower[12'd447] = 8'd120;
vramDataLower[12'd448] = 8'd207;
vramDataLower[12'd449] = 8'd120;
vramDataLower[12'd450] = 8'd31;
vramDataLower[12'd451] = 8'd120;
vramDataLower[12'd452] = 8'd30;
vramDataLower[12'd453] = 8'd120;
vramDataLower[12'd454] = 8'd183;
vramDataLower[12'd455] = 8'd120;
vramDataLower[12'd456] = 8'd198;
vramDataLower[12'd457] = 8'd120;
vramDataLower[12'd458] = 8'd135;
vramDataLower[12'd459] = 8'd135;
vramDataLower[12'd460] = 8'd52;
vramDataLower[12'd461] = 8'd87;
vramDataLower[12'd462] = 8'd70;
vramDataLower[12'd463] = 8'd87;
vramDataLower[12'd464] = 8'd39;
vramDataLower[12'd465] = 8'd247;
vramDataLower[12'd466] = 8'd16;
vramDataLower[12'd467] = 8'd247;
vramDataLower[12'd468] = 8'd146;
vramDataLower[12'd469] = 8'd119;
vramDataLower[12'd470] = 8'd255;
vramDataLower[12'd471] = 8'd199;
vramDataLower[12'd472] = 8'd210;
vramDataLower[12'd473] = 8'd55;
vramDataLower[12'd474] = 8'd210;
vramDataLower[12'd475] = 8'd55;
vramDataLower[12'd476] = 8'd164;
vramDataLower[12'd477] = 8'd152;
vramDataLower[12'd478] = 8'd16;
vramDataLower[12'd479] = 8'd135;
vramDataLower[12'd480] = 8'd210;
vramDataLower[12'd481] = 8'd55;
vramDataLower[12'd482] = 8'd202;
vramDataLower[12'd483] = 8'd183;
vramDataLower[12'd484] = 8'd202;
vramDataLower[12'd485] = 8'd183;
vramDataLower[12'd486] = 8'd202;
vramDataLower[12'd487] = 8'd183;
vramDataLower[12'd488] = 8'd202;
vramDataLower[12'd489] = 8'd183;
vramDataLower[12'd490] = 8'd202;
vramDataLower[12'd491] = 8'd183;
vramDataLower[12'd492] = 8'd202;
vramDataLower[12'd493] = 8'd183;
vramDataLower[12'd494] = 8'd202;
vramDataLower[12'd495] = 8'd183;
vramDataLower[12'd496] = 8'd202;
vramDataLower[12'd497] = 8'd183;
vramDataLower[12'd498] = 8'd202;
vramDataLower[12'd499] = 8'd183;
vramDataLower[12'd500] = 8'd31;
vramDataLower[12'd501] = 8'd183;
vramDataLower[12'd502] = 8'd31;
vramDataLower[12'd503] = 8'd183;
vramDataLower[12'd504] = 8'd48;
vramDataLower[12'd505] = 8'd183;
vramDataLower[12'd506] = 8'd37;
vramDataLower[12'd507] = 8'd183;
vramDataLower[12'd508] = 8'd202;
vramDataLower[12'd509] = 8'd183;
vramDataLower[12'd510] = 8'd202;
vramDataLower[12'd511] = 8'd183;
vramDataLower[12'd512] = 8'd202;
vramDataLower[12'd513] = 8'd183;
vramDataLower[12'd514] = 8'd202;
vramDataLower[12'd515] = 8'd183;
vramDataLower[12'd516] = 8'd202;
vramDataLower[12'd517] = 8'd183;
vramDataLower[12'd518] = 8'd202;
vramDataLower[12'd519] = 8'd183;
vramDataLower[12'd520] = 8'd16;
vramDataLower[12'd521] = 8'd183;
vramDataLower[12'd522] = 8'd16;
vramDataLower[12'd523] = 8'd247;
vramDataLower[12'd524] = 8'd16;
vramDataLower[12'd525] = 8'd183;
vramDataLower[12'd526] = 8'd181;
vramDataLower[12'd527] = 8'd135;
vramDataLower[12'd528] = 8'd188;
vramDataLower[12'd529] = 8'd135;
vramDataLower[12'd530] = 8'd252;
vramDataLower[12'd531] = 8'd135;
vramDataLower[12'd532] = 8'd248;
vramDataLower[12'd533] = 8'd55;
vramDataLower[12'd534] = 8'd249;
vramDataLower[12'd535] = 8'd247;
vramDataLower[12'd536] = 8'd40;
vramDataLower[12'd537] = 8'd119;
vramDataLower[12'd538] = 8'd95;
vramDataLower[12'd539] = 8'd55;
vramDataLower[12'd540] = 8'd214;
vramDataLower[12'd541] = 8'd55;
vramDataLower[12'd542] = 8'd183;
vramDataLower[12'd543] = 8'd55;
vramDataLower[12'd544] = 8'd44;
vramDataLower[12'd545] = 8'd87;
vramDataLower[12'd546] = 8'd7;
vramDataLower[12'd547] = 8'd87;
vramDataLower[12'd548] = 8'd97;
vramDataLower[12'd549] = 8'd119;
vramDataLower[12'd550] = 8'd95;
vramDataLower[12'd551] = 8'd55;
vramDataLower[12'd552] = 8'd39;
vramDataLower[12'd553] = 8'd247;
vramDataLower[12'd554] = 8'd32;
vramDataLower[12'd555] = 8'd183;
vramDataLower[12'd556] = 8'd16;
vramDataLower[12'd557] = 8'd247;
vramDataLower[12'd558] = 8'd170;
vramDataLower[12'd559] = 8'd247;
vramDataLower[12'd560] = 8'd249;
vramDataLower[12'd561] = 8'd87;
vramDataLower[12'd562] = 8'd217;
vramDataLower[12'd563] = 8'd247;
vramDataLower[12'd564] = 8'd209;
vramDataLower[12'd565] = 8'd247;
vramDataLower[12'd566] = 8'd106;
vramDataLower[12'd567] = 8'd247;
vramDataLower[12'd568] = 8'd31;
vramDataLower[12'd569] = 8'd247;
vramDataLower[12'd570] = 8'd94;
vramDataLower[12'd571] = 8'd55;
vramDataLower[12'd572] = 8'd17;
vramDataLower[12'd573] = 8'd247;
vramDataLower[12'd574] = 8'd17;
vramDataLower[12'd575] = 8'd247;
vramDataLower[12'd576] = 8'd202;
vramDataLower[12'd577] = 8'd247;
vramDataLower[12'd578] = 8'd7;
vramDataLower[12'd579] = 8'd247;
vramDataLower[12'd580] = 8'd117;
vramDataLower[12'd581] = 8'd247;
vramDataLower[12'd582] = 8'd200;
vramDataLower[12'd583] = 8'd135;
vramDataLower[12'd584] = 8'd220;
vramDataLower[12'd585] = 8'd120;
vramDataLower[12'd586] = 8'd223;
vramDataLower[12'd587] = 8'd135;
vramDataLower[12'd588] = 8'd95;
vramDataLower[12'd589] = 8'd135;
vramDataLower[12'd590] = 8'd210;
vramDataLower[12'd591] = 8'd135;
vramDataLower[12'd592] = 8'd188;
vramDataLower[12'd593] = 8'd120;
vramDataLower[12'd594] = 8'd150;
vramDataLower[12'd595] = 8'd152;
vramDataLower[12'd596] = 8'd16;
vramDataLower[12'd597] = 8'd152;
vramDataLower[12'd598] = 8'd183;
vramDataLower[12'd599] = 8'd136;
vramDataLower[12'd600] = 8'd46;
vramDataLower[12'd601] = 8'd152;
vramDataLower[12'd602] = 8'd214;
vramDataLower[12'd603] = 8'd152;
vramDataLower[12'd604] = 8'd200;
vramDataLower[12'd605] = 8'd120;
vramDataLower[12'd606] = 8'd80;
vramDataLower[12'd607] = 8'd120;
vramDataLower[12'd608] = 8'd55;
vramDataLower[12'd609] = 8'd120;
vramDataLower[12'd610] = 8'd126;
vramDataLower[12'd611] = 8'd120;
vramDataLower[12'd612] = 8'd202;
vramDataLower[12'd613] = 8'd120;
vramDataLower[12'd614] = 8'd31;
vramDataLower[12'd615] = 8'd120;
vramDataLower[12'd616] = 8'd202;
vramDataLower[12'd617] = 8'd135;
vramDataLower[12'd618] = 8'd202;
vramDataLower[12'd619] = 8'd135;
vramDataLower[12'd620] = 8'd16;
vramDataLower[12'd621] = 8'd87;
vramDataLower[12'd622] = 8'd31;
vramDataLower[12'd623] = 8'd247;
vramDataLower[12'd624] = 8'd230;
vramDataLower[12'd625] = 8'd247;
vramDataLower[12'd626] = 8'd156;
vramDataLower[12'd627] = 8'd247;
vramDataLower[12'd628] = 8'd65;
vramDataLower[12'd629] = 8'd119;
vramDataLower[12'd630] = 8'd214;
vramDataLower[12'd631] = 8'd55;
vramDataLower[12'd632] = 8'd210;
vramDataLower[12'd633] = 8'd55;
vramDataLower[12'd634] = 8'd214;
vramDataLower[12'd635] = 8'd135;
vramDataLower[12'd636] = 8'd164;
vramDataLower[12'd637] = 8'd120;
vramDataLower[12'd638] = 8'd16;
vramDataLower[12'd639] = 8'd127;
vramDataLower[12'd640] = 8'd16;
vramDataLower[12'd641] = 8'd8;
vramDataLower[12'd642] = 8'd230;
vramDataLower[12'd643] = 8'd135;
vramDataLower[12'd644] = 8'd31;
vramDataLower[12'd645] = 8'd247;
vramDataLower[12'd646] = 8'd31;
vramDataLower[12'd647] = 8'd247;
vramDataLower[12'd648] = 8'd31;
vramDataLower[12'd649] = 8'd247;
vramDataLower[12'd650] = 8'd30;
vramDataLower[12'd651] = 8'd247;
vramDataLower[12'd652] = 8'd30;
vramDataLower[12'd653] = 8'd247;
vramDataLower[12'd654] = 8'd30;
vramDataLower[12'd655] = 8'd247;
vramDataLower[12'd656] = 8'd30;
vramDataLower[12'd657] = 8'd247;
vramDataLower[12'd658] = 8'd30;
vramDataLower[12'd659] = 8'd247;
vramDataLower[12'd660] = 8'd30;
vramDataLower[12'd661] = 8'd247;
vramDataLower[12'd662] = 8'd210;
vramDataLower[12'd663] = 8'd247;
vramDataLower[12'd664] = 8'd183;
vramDataLower[12'd665] = 8'd247;
vramDataLower[12'd666] = 8'd183;
vramDataLower[12'd667] = 8'd247;
vramDataLower[12'd668] = 8'd252;
vramDataLower[12'd669] = 8'd55;
vramDataLower[12'd670] = 8'd252;
vramDataLower[12'd671] = 8'd55;
vramDataLower[12'd672] = 8'd252;
vramDataLower[12'd673] = 8'd55;
vramDataLower[12'd674] = 8'd252;
vramDataLower[12'd675] = 8'd55;
vramDataLower[12'd676] = 8'd166;
vramDataLower[12'd677] = 8'd55;
vramDataLower[12'd678] = 8'd126;
vramDataLower[12'd679] = 8'd55;
vramDataLower[12'd680] = 8'd39;
vramDataLower[12'd681] = 8'd55;
vramDataLower[12'd682] = 8'd94;
vramDataLower[12'd683] = 8'd247;
vramDataLower[12'd684] = 8'd237;
vramDataLower[12'd685] = 8'd119;
vramDataLower[12'd686] = 8'd210;
vramDataLower[12'd687] = 8'd55;
vramDataLower[12'd688] = 8'd230;
vramDataLower[12'd689] = 8'd135;
vramDataLower[12'd690] = 8'd249;
vramDataLower[12'd691] = 8'd55;
vramDataLower[12'd692] = 8'd213;
vramDataLower[12'd693] = 8'd55;
vramDataLower[12'd694] = 8'd230;
vramDataLower[12'd695] = 8'd135;
vramDataLower[12'd696] = 8'd198;
vramDataLower[12'd697] = 8'd135;
vramDataLower[12'd698] = 8'd198;
vramDataLower[12'd699] = 8'd135;
vramDataLower[12'd700] = 8'd16;
vramDataLower[12'd701] = 8'd135;
vramDataLower[12'd702] = 8'd230;
vramDataLower[12'd703] = 8'd135;
vramDataLower[12'd704] = 8'd230;
vramDataLower[12'd705] = 8'd135;
vramDataLower[12'd706] = 8'd19;
vramDataLower[12'd707] = 8'd135;
vramDataLower[12'd708] = 8'd17;
vramDataLower[12'd709] = 8'd55;
vramDataLower[12'd710] = 8'd96;
vramDataLower[12'd711] = 8'd55;
vramDataLower[12'd712] = 8'd0;
vramDataLower[12'd713] = 8'd71;
vramDataLower[12'd714] = 8'd44;
vramDataLower[12'd715] = 8'd135;
vramDataLower[12'd716] = 8'd96;
vramDataLower[12'd717] = 8'd247;
vramDataLower[12'd718] = 8'd251;
vramDataLower[12'd719] = 8'd247;
vramDataLower[12'd720] = 8'd212;
vramDataLower[12'd721] = 8'd247;
vramDataLower[12'd722] = 8'd44;
vramDataLower[12'd723] = 8'd247;
vramDataLower[12'd724] = 8'd249;
vramDataLower[12'd725] = 8'd55;
vramDataLower[12'd726] = 8'd7;
vramDataLower[12'd727] = 8'd55;
vramDataLower[12'd728] = 8'd250;
vramDataLower[12'd729] = 8'd247;
vramDataLower[12'd730] = 8'd166;
vramDataLower[12'd731] = 8'd55;
vramDataLower[12'd732] = 8'd135;
vramDataLower[12'd733] = 8'd247;
vramDataLower[12'd734] = 8'd44;
vramDataLower[12'd735] = 8'd103;
vramDataLower[12'd736] = 8'd192;
vramDataLower[12'd737] = 8'd135;
vramDataLower[12'd738] = 8'd17;
vramDataLower[12'd739] = 8'd135;
vramDataLower[12'd740] = 8'd214;
vramDataLower[12'd741] = 8'd135;
vramDataLower[12'd742] = 8'd16;
vramDataLower[12'd743] = 8'd135;
vramDataLower[12'd744] = 8'd183;
vramDataLower[12'd745] = 8'd135;
vramDataLower[12'd746] = 8'd214;
vramDataLower[12'd747] = 8'd135;
vramDataLower[12'd748] = 8'd148;
vramDataLower[12'd749] = 8'd120;
vramDataLower[12'd750] = 8'd16;
vramDataLower[12'd751] = 8'd120;
vramDataLower[12'd752] = 8'd135;
vramDataLower[12'd753] = 8'd120;
vramDataLower[12'd754] = 8'd230;
vramDataLower[12'd755] = 8'd120;
vramDataLower[12'd756] = 8'd76;
vramDataLower[12'd757] = 8'd120;
vramDataLower[12'd758] = 8'd95;
vramDataLower[12'd759] = 8'd120;
vramDataLower[12'd760] = 8'd31;
vramDataLower[12'd761] = 8'd152;
vramDataLower[12'd762] = 8'd102;
vramDataLower[12'd763] = 8'd120;
vramDataLower[12'd764] = 8'd9;
vramDataLower[12'd765] = 8'd120;
vramDataLower[12'd766] = 8'd202;
vramDataLower[12'd767] = 8'd120;
vramDataLower[12'd768] = 8'd31;
vramDataLower[12'd769] = 8'd120;
vramDataLower[12'd770] = 8'd202;
vramDataLower[12'd771] = 8'd120;
vramDataLower[12'd772] = 8'd164;
vramDataLower[12'd773] = 8'd135;
vramDataLower[12'd774] = 8'd230;
vramDataLower[12'd775] = 8'd135;
vramDataLower[12'd776] = 8'd126;
vramDataLower[12'd777] = 8'd135;
vramDataLower[12'd778] = 8'd167;
vramDataLower[12'd779] = 8'd135;
vramDataLower[12'd780] = 8'd46;
vramDataLower[12'd781] = 8'd135;
vramDataLower[12'd782] = 8'd214;
vramDataLower[12'd783] = 8'd247;
vramDataLower[12'd784] = 8'd253;
vramDataLower[12'd785] = 8'd247;
vramDataLower[12'd786] = 8'd96;
vramDataLower[12'd787] = 8'd247;
vramDataLower[12'd788] = 8'd214;
vramDataLower[12'd789] = 8'd55;
vramDataLower[12'd790] = 8'd210;
vramDataLower[12'd791] = 8'd55;
vramDataLower[12'd792] = 8'd210;
vramDataLower[12'd793] = 8'd55;
vramDataLower[12'd794] = 8'd16;
vramDataLower[12'd795] = 8'd120;
vramDataLower[12'd796] = 8'd221;
vramDataLower[12'd797] = 8'd135;
vramDataLower[12'd798] = 8'd85;
vramDataLower[12'd799] = 8'd127;
vramDataLower[12'd800] = 8'd202;
vramDataLower[12'd801] = 8'd8;
vramDataLower[12'd802] = 8'd16;
vramDataLower[12'd803] = 8'd8;
vramDataLower[12'd804] = 8'd16;
vramDataLower[12'd805] = 8'd135;
vramDataLower[12'd806] = 8'd16;
vramDataLower[12'd807] = 8'd103;
vramDataLower[12'd808] = 8'd16;
vramDataLower[12'd809] = 8'd103;
vramDataLower[12'd810] = 8'd30;
vramDataLower[12'd811] = 8'd103;
vramDataLower[12'd812] = 8'd16;
vramDataLower[12'd813] = 8'd103;
vramDataLower[12'd814] = 8'd164;
vramDataLower[12'd815] = 8'd103;
vramDataLower[12'd816] = 8'd209;
vramDataLower[12'd817] = 8'd231;
vramDataLower[12'd818] = 8'd210;
vramDataLower[12'd819] = 8'd247;
vramDataLower[12'd820] = 8'd210;
vramDataLower[12'd821] = 8'd247;
vramDataLower[12'd822] = 8'd210;
vramDataLower[12'd823] = 8'd247;
vramDataLower[12'd824] = 8'd210;
vramDataLower[12'd825] = 8'd247;
vramDataLower[12'd826] = 8'd30;
vramDataLower[12'd827] = 8'd247;
vramDataLower[12'd828] = 8'd95;
vramDataLower[12'd829] = 8'd247;
vramDataLower[12'd830] = 8'd250;
vramDataLower[12'd831] = 8'd247;
vramDataLower[12'd832] = 8'd94;
vramDataLower[12'd833] = 8'd247;
vramDataLower[12'd834] = 8'd94;
vramDataLower[12'd835] = 8'd247;
vramDataLower[12'd836] = 8'd189;
vramDataLower[12'd837] = 8'd119;
vramDataLower[12'd838] = 8'd95;
vramDataLower[12'd839] = 8'd55;
vramDataLower[12'd840] = 8'd210;
vramDataLower[12'd841] = 8'd55;
vramDataLower[12'd842] = 8'd214;
vramDataLower[12'd843] = 8'd135;
vramDataLower[12'd844] = 8'd210;
vramDataLower[12'd845] = 8'd135;
vramDataLower[12'd846] = 8'd198;
vramDataLower[12'd847] = 8'd135;
vramDataLower[12'd848] = 8'd16;
vramDataLower[12'd849] = 8'd135;
vramDataLower[12'd850] = 8'd16;
vramDataLower[12'd851] = 8'd135;
vramDataLower[12'd852] = 8'd80;
vramDataLower[12'd853] = 8'd120;
vramDataLower[12'd854] = 8'd202;
vramDataLower[12'd855] = 8'd120;
vramDataLower[12'd856] = 8'd16;
vramDataLower[12'd857] = 8'd135;
vramDataLower[12'd858] = 8'd159;
vramDataLower[12'd859] = 8'd135;
vramDataLower[12'd860] = 8'd16;
vramDataLower[12'd861] = 8'd120;
vramDataLower[12'd862] = 8'd135;
vramDataLower[12'd863] = 8'd135;
vramDataLower[12'd864] = 8'd37;
vramDataLower[12'd865] = 8'd135;
vramDataLower[12'd866] = 8'd17;
vramDataLower[12'd867] = 8'd135;
vramDataLower[12'd868] = 8'd53;
vramDataLower[12'd869] = 8'd119;
vramDataLower[12'd870] = 8'd179;
vramDataLower[12'd871] = 8'd87;
vramDataLower[12'd872] = 8'd95;
vramDataLower[12'd873] = 8'd87;
vramDataLower[12'd874] = 8'd96;
vramDataLower[12'd875] = 8'd135;
vramDataLower[12'd876] = 8'd214;
vramDataLower[12'd877] = 8'd247;
vramDataLower[12'd878] = 8'd183;
vramDataLower[12'd879] = 8'd103;
vramDataLower[12'd880] = 8'd126;
vramDataLower[12'd881] = 8'd247;
vramDataLower[12'd882] = 8'd94;
vramDataLower[12'd883] = 8'd247;
vramDataLower[12'd884] = 8'd226;
vramDataLower[12'd885] = 8'd247;
vramDataLower[12'd886] = 8'd39;
vramDataLower[12'd887] = 8'd247;
vramDataLower[12'd888] = 8'd152;
vramDataLower[12'd889] = 8'd119;
vramDataLower[12'd890] = 8'd39;
vramDataLower[12'd891] = 8'd247;
vramDataLower[12'd892] = 8'd44;
vramDataLower[12'd893] = 8'd135;
vramDataLower[12'd894] = 8'd189;
vramDataLower[12'd895] = 8'd103;
vramDataLower[12'd896] = 8'd95;
vramDataLower[12'd897] = 8'd135;
vramDataLower[12'd898] = 8'd90;
vramDataLower[12'd899] = 8'd135;
vramDataLower[12'd900] = 8'd202;
vramDataLower[12'd901] = 8'd135;
vramDataLower[12'd902] = 8'd17;
vramDataLower[12'd903] = 8'd120;
vramDataLower[12'd904] = 8'd85;
vramDataLower[12'd905] = 8'd135;
vramDataLower[12'd906] = 8'd16;
vramDataLower[12'd907] = 8'd120;
vramDataLower[12'd908] = 8'd210;
vramDataLower[12'd909] = 8'd120;
vramDataLower[12'd910] = 8'd188;
vramDataLower[12'd911] = 8'd120;
vramDataLower[12'd912] = 8'd202;
vramDataLower[12'd913] = 8'd120;
vramDataLower[12'd914] = 8'd253;
vramDataLower[12'd915] = 8'd120;
vramDataLower[12'd916] = 8'd198;
vramDataLower[12'd917] = 8'd120;
vramDataLower[12'd918] = 8'd198;
vramDataLower[12'd919] = 8'd120;
vramDataLower[12'd920] = 8'd230;
vramDataLower[12'd921] = 8'd120;
vramDataLower[12'd922] = 8'd16;
vramDataLower[12'd923] = 8'd120;
vramDataLower[12'd924] = 8'd9;
vramDataLower[12'd925] = 8'd120;
vramDataLower[12'd926] = 8'd31;
vramDataLower[12'd927] = 8'd120;
vramDataLower[12'd928] = 8'd37;
vramDataLower[12'd929] = 8'd120;
vramDataLower[12'd930] = 8'd85;
vramDataLower[12'd931] = 8'd120;
vramDataLower[12'd932] = 8'd37;
vramDataLower[12'd933] = 8'd120;
vramDataLower[12'd934] = 8'd210;
vramDataLower[12'd935] = 8'd135;
vramDataLower[12'd936] = 8'd183;
vramDataLower[12'd937] = 8'd135;
vramDataLower[12'd938] = 8'd17;
vramDataLower[12'd939] = 8'd135;
vramDataLower[12'd940] = 8'd29;
vramDataLower[12'd941] = 8'd247;
vramDataLower[12'd942] = 8'd229;
vramDataLower[12'd943] = 8'd247;
vramDataLower[12'd944] = 8'd46;
vramDataLower[12'd945] = 8'd247;
vramDataLower[12'd946] = 8'd210;
vramDataLower[12'd947] = 8'd55;
vramDataLower[12'd948] = 8'd210;
vramDataLower[12'd949] = 8'd135;
vramDataLower[12'd950] = 8'd210;
vramDataLower[12'd951] = 8'd135;
vramDataLower[12'd952] = 8'd210;
vramDataLower[12'd953] = 8'd135;
vramDataLower[12'd954] = 8'd70;
vramDataLower[12'd955] = 8'd120;
vramDataLower[12'd956] = 8'd16;
vramDataLower[12'd957] = 8'd135;
vramDataLower[12'd958] = 8'd80;
vramDataLower[12'd959] = 8'd123;
vramDataLower[12'd960] = 8'd210;
vramDataLower[12'd961] = 8'd8;
vramDataLower[12'd962] = 8'd65;
vramDataLower[12'd963] = 8'd136;
vramDataLower[12'd964] = 8'd135;
vramDataLower[12'd965] = 8'd135;
vramDataLower[12'd966] = 8'd210;
vramDataLower[12'd967] = 8'd103;
vramDataLower[12'd968] = 8'd210;
vramDataLower[12'd969] = 8'd103;
vramDataLower[12'd970] = 8'd210;
vramDataLower[12'd971] = 8'd103;
vramDataLower[12'd972] = 8'd210;
vramDataLower[12'd973] = 8'd103;
vramDataLower[12'd974] = 8'd183;
vramDataLower[12'd975] = 8'd103;
vramDataLower[12'd976] = 8'd202;
vramDataLower[12'd977] = 8'd231;
vramDataLower[12'd978] = 8'd30;
vramDataLower[12'd979] = 8'd247;
vramDataLower[12'd980] = 8'd30;
vramDataLower[12'd981] = 8'd247;
vramDataLower[12'd982] = 8'd30;
vramDataLower[12'd983] = 8'd247;
vramDataLower[12'd984] = 8'd16;
vramDataLower[12'd985] = 8'd247;
vramDataLower[12'd986] = 8'd16;
vramDataLower[12'd987] = 8'd247;
vramDataLower[12'd988] = 8'd45;
vramDataLower[12'd989] = 8'd247;
vramDataLower[12'd990] = 8'd95;
vramDataLower[12'd991] = 8'd135;
vramDataLower[12'd992] = 8'd183;
vramDataLower[12'd993] = 8'd135;
vramDataLower[12'd994] = 8'd209;
vramDataLower[12'd995] = 8'd135;
vramDataLower[12'd996] = 8'd210;
vramDataLower[12'd997] = 8'd135;
vramDataLower[12'd998] = 8'd202;
vramDataLower[12'd999] = 8'd120;
vramDataLower[12'd1000] = 8'd80;
vramDataLower[12'd1001] = 8'd120;
vramDataLower[12'd1002] = 8'd202;
vramDataLower[12'd1003] = 8'd152;
vramDataLower[12'd1004] = 8'd198;
vramDataLower[12'd1005] = 8'd152;
vramDataLower[12'd1006] = 8'd200;
vramDataLower[12'd1007] = 8'd120;
vramDataLower[12'd1008] = 8'd181;
vramDataLower[12'd1009] = 8'd120;
vramDataLower[12'd1010] = 8'd85;
vramDataLower[12'd1011] = 8'd120;
vramDataLower[12'd1012] = 8'd181;
vramDataLower[12'd1013] = 8'd135;
vramDataLower[12'd1014] = 8'd135;
vramDataLower[12'd1015] = 8'd120;
vramDataLower[12'd1016] = 8'd208;
vramDataLower[12'd1017] = 8'd120;
vramDataLower[12'd1018] = 8'd188;
vramDataLower[12'd1019] = 8'd120;
vramDataLower[12'd1020] = 8'd30;
vramDataLower[12'd1021] = 8'd120;
vramDataLower[12'd1022] = 8'd164;
vramDataLower[12'd1023] = 8'd120;
vramDataLower[12'd1024] = 8'd148;
vramDataLower[12'd1025] = 8'd135;
vramDataLower[12'd1026] = 8'd17;
vramDataLower[12'd1027] = 8'd135;
vramDataLower[12'd1028] = 8'd209;
vramDataLower[12'd1029] = 8'd55;
vramDataLower[12'd1030] = 8'd198;
vramDataLower[12'd1031] = 8'd135;
vramDataLower[12'd1032] = 8'd16;
vramDataLower[12'd1033] = 8'd135;
vramDataLower[12'd1034] = 8'd95;
vramDataLower[12'd1035] = 8'd135;
vramDataLower[12'd1036] = 8'd12;
vramDataLower[12'd1037] = 8'd119;
vramDataLower[12'd1038] = 8'd180;
vramDataLower[12'd1039] = 8'd87;
vramDataLower[12'd1040] = 8'd183;
vramDataLower[12'd1041] = 8'd103;
vramDataLower[12'd1042] = 8'd7;
vramDataLower[12'd1043] = 8'd135;
vramDataLower[12'd1044] = 8'd213;
vramDataLower[12'd1045] = 8'd55;
vramDataLower[12'd1046] = 8'd210;
vramDataLower[12'd1047] = 8'd135;
vramDataLower[12'd1048] = 8'd85;
vramDataLower[12'd1049] = 8'd120;
vramDataLower[12'd1050] = 8'd248;
vramDataLower[12'd1051] = 8'd120;
vramDataLower[12'd1052] = 8'd198;
vramDataLower[12'd1053] = 8'd120;
vramDataLower[12'd1054] = 8'd210;
vramDataLower[12'd1055] = 8'd135;
vramDataLower[12'd1056] = 8'd109;
vramDataLower[12'd1057] = 8'd135;
vramDataLower[12'd1058] = 8'd16;
vramDataLower[12'd1059] = 8'd135;
vramDataLower[12'd1060] = 8'd210;
vramDataLower[12'd1061] = 8'd135;
vramDataLower[12'd1062] = 8'd181;
vramDataLower[12'd1063] = 8'd135;
vramDataLower[12'd1064] = 8'd210;
vramDataLower[12'd1065] = 8'd135;
vramDataLower[12'd1066] = 8'd85;
vramDataLower[12'd1067] = 8'd135;
vramDataLower[12'd1068] = 8'd90;
vramDataLower[12'd1069] = 8'd120;
vramDataLower[12'd1070] = 8'd210;
vramDataLower[12'd1071] = 8'd120;
vramDataLower[12'd1072] = 8'd16;
vramDataLower[12'd1073] = 8'd120;
vramDataLower[12'd1074] = 8'd31;
vramDataLower[12'd1075] = 8'd120;
vramDataLower[12'd1076] = 8'd30;
vramDataLower[12'd1077] = 8'd120;
vramDataLower[12'd1078] = 8'd164;
vramDataLower[12'd1079] = 8'd120;
vramDataLower[12'd1080] = 8'd16;
vramDataLower[12'd1081] = 8'd120;
vramDataLower[12'd1082] = 8'd213;
vramDataLower[12'd1083] = 8'd120;
vramDataLower[12'd1084] = 8'd210;
vramDataLower[12'd1085] = 8'd120;
vramDataLower[12'd1086] = 8'd16;
vramDataLower[12'd1087] = 8'd120;
vramDataLower[12'd1088] = 8'd202;
vramDataLower[12'd1089] = 8'd135;
vramDataLower[12'd1090] = 8'd202;
vramDataLower[12'd1091] = 8'd135;
vramDataLower[12'd1092] = 8'd248;
vramDataLower[12'd1093] = 8'd135;
vramDataLower[12'd1094] = 8'd126;
vramDataLower[12'd1095] = 8'd135;
vramDataLower[12'd1096] = 8'd248;
vramDataLower[12'd1097] = 8'd135;
vramDataLower[12'd1098] = 8'd55;
vramDataLower[12'd1099] = 8'd135;
vramDataLower[12'd1100] = 8'd37;
vramDataLower[12'd1101] = 8'd55;
vramDataLower[12'd1102] = 8'd31;
vramDataLower[12'd1103] = 8'd135;
vramDataLower[12'd1104] = 8'd34;
vramDataLower[12'd1105] = 8'd247;
vramDataLower[12'd1106] = 8'd200;
vramDataLower[12'd1107] = 8'd55;
vramDataLower[12'd1108] = 8'd202;
vramDataLower[12'd1109] = 8'd55;
vramDataLower[12'd1110] = 8'd83;
vramDataLower[12'd1111] = 8'd135;
vramDataLower[12'd1112] = 8'd80;
vramDataLower[12'd1113] = 8'd120;
vramDataLower[12'd1114] = 8'd210;
vramDataLower[12'd1115] = 8'd120;
vramDataLower[12'd1116] = 8'd210;
vramDataLower[12'd1117] = 8'd55;
vramDataLower[12'd1118] = 8'd202;
vramDataLower[12'd1119] = 8'd179;
vramDataLower[12'd1120] = 8'd16;
vramDataLower[12'd1121] = 8'd24;
vramDataLower[12'd1122] = 8'd214;
vramDataLower[12'd1123] = 8'd120;
vramDataLower[12'd1124] = 8'd220;
vramDataLower[12'd1125] = 8'd120;
vramDataLower[12'd1126] = 8'd220;
vramDataLower[12'd1127] = 8'd120;
vramDataLower[12'd1128] = 8'd223;
vramDataLower[12'd1129] = 8'd135;
vramDataLower[12'd1130] = 8'd223;
vramDataLower[12'd1131] = 8'd135;
vramDataLower[12'd1132] = 8'd223;
vramDataLower[12'd1133] = 8'd135;
vramDataLower[12'd1134] = 8'd220;
vramDataLower[12'd1135] = 8'd120;
vramDataLower[12'd1136] = 8'd223;
vramDataLower[12'd1137] = 8'd135;
vramDataLower[12'd1138] = 8'd31;
vramDataLower[12'd1139] = 8'd135;
vramDataLower[12'd1140] = 8'd31;
vramDataLower[12'd1141] = 8'd135;
vramDataLower[12'd1142] = 8'd31;
vramDataLower[12'd1143] = 8'd135;
vramDataLower[12'd1144] = 8'd31;
vramDataLower[12'd1145] = 8'd135;
vramDataLower[12'd1146] = 8'd30;
vramDataLower[12'd1147] = 8'd135;
vramDataLower[12'd1148] = 8'd210;
vramDataLower[12'd1149] = 8'd135;
vramDataLower[12'd1150] = 8'd202;
vramDataLower[12'd1151] = 8'd120;
vramDataLower[12'd1152] = 8'd248;
vramDataLower[12'd1153] = 8'd120;
vramDataLower[12'd1154] = 8'd94;
vramDataLower[12'd1155] = 8'd120;
vramDataLower[12'd1156] = 8'd211;
vramDataLower[12'd1157] = 8'd120;
vramDataLower[12'd1158] = 8'd16;
vramDataLower[12'd1159] = 8'd120;
vramDataLower[12'd1160] = 8'd94;
vramDataLower[12'd1161] = 8'd152;
vramDataLower[12'd1162] = 8'd94;
vramDataLower[12'd1163] = 8'd8;
vramDataLower[12'd1164] = 8'd212;
vramDataLower[12'd1165] = 8'd152;
vramDataLower[12'd1166] = 8'd181;
vramDataLower[12'd1167] = 8'd152;
vramDataLower[12'd1168] = 8'd202;
vramDataLower[12'd1169] = 8'd152;
vramDataLower[12'd1170] = 8'd166;
vramDataLower[12'd1171] = 8'd120;
vramDataLower[12'd1172] = 8'd210;
vramDataLower[12'd1173] = 8'd120;
vramDataLower[12'd1174] = 8'd85;
vramDataLower[12'd1175] = 8'd120;
vramDataLower[12'd1176] = 8'd148;
vramDataLower[12'd1177] = 8'd120;
vramDataLower[12'd1178] = 8'd230;
vramDataLower[12'd1179] = 8'd120;
vramDataLower[12'd1180] = 8'd164;
vramDataLower[12'd1181] = 8'd152;
vramDataLower[12'd1182] = 8'd194;
vramDataLower[12'd1183] = 8'd120;
vramDataLower[12'd1184] = 8'd80;
vramDataLower[12'd1185] = 8'd135;
vramDataLower[12'd1186] = 8'd181;
vramDataLower[12'd1187] = 8'd135;
vramDataLower[12'd1188] = 8'd16;
vramDataLower[12'd1189] = 8'd135;
vramDataLower[12'd1190] = 8'd31;
vramDataLower[12'd1191] = 8'd135;
vramDataLower[12'd1192] = 8'd164;
vramDataLower[12'd1193] = 8'd135;
vramDataLower[12'd1194] = 8'd218;
vramDataLower[12'd1195] = 8'd135;
vramDataLower[12'd1196] = 8'd184;
vramDataLower[12'd1197] = 8'd135;
vramDataLower[12'd1198] = 8'd95;
vramDataLower[12'd1199] = 8'd87;
vramDataLower[12'd1200] = 8'd95;
vramDataLower[12'd1201] = 8'd135;
vramDataLower[12'd1202] = 8'd202;
vramDataLower[12'd1203] = 8'd120;
vramDataLower[12'd1204] = 8'd80;
vramDataLower[12'd1205] = 8'd120;
vramDataLower[12'd1206] = 8'd252;
vramDataLower[12'd1207] = 8'd120;
vramDataLower[12'd1208] = 8'd202;
vramDataLower[12'd1209] = 8'd120;
vramDataLower[12'd1210] = 8'd85;
vramDataLower[12'd1211] = 8'd120;
vramDataLower[12'd1212] = 8'd150;
vramDataLower[12'd1213] = 8'd120;
vramDataLower[12'd1214] = 8'd172;
vramDataLower[12'd1215] = 8'd135;
vramDataLower[12'd1216] = 8'd164;
vramDataLower[12'd1217] = 8'd135;
vramDataLower[12'd1218] = 8'd202;
vramDataLower[12'd1219] = 8'd120;
vramDataLower[12'd1220] = 8'd181;
vramDataLower[12'd1221] = 8'd120;
vramDataLower[12'd1222] = 8'd210;
vramDataLower[12'd1223] = 8'd120;
vramDataLower[12'd1224] = 8'd85;
vramDataLower[12'd1225] = 8'd120;
vramDataLower[12'd1226] = 8'd230;
vramDataLower[12'd1227] = 8'd135;
vramDataLower[12'd1228] = 8'd171;
vramDataLower[12'd1229] = 8'd135;
vramDataLower[12'd1230] = 8'd198;
vramDataLower[12'd1231] = 8'd135;
vramDataLower[12'd1232] = 8'd197;
vramDataLower[12'd1233] = 8'd135;
vramDataLower[12'd1234] = 8'd230;
vramDataLower[12'd1235] = 8'd120;
vramDataLower[12'd1236] = 8'd210;
vramDataLower[12'd1237] = 8'd120;
vramDataLower[12'd1238] = 8'd31;
vramDataLower[12'd1239] = 8'd120;
vramDataLower[12'd1240] = 8'd135;
vramDataLower[12'd1241] = 8'd120;
vramDataLower[12'd1242] = 8'd31;
vramDataLower[12'd1243] = 8'd120;
vramDataLower[12'd1244] = 8'd31;
vramDataLower[12'd1245] = 8'd120;
vramDataLower[12'd1246] = 8'd16;
vramDataLower[12'd1247] = 8'd135;
vramDataLower[12'd1248] = 8'd214;
vramDataLower[12'd1249] = 8'd135;
vramDataLower[12'd1250] = 8'd30;
vramDataLower[12'd1251] = 8'd87;
vramDataLower[12'd1252] = 8'd16;
vramDataLower[12'd1253] = 8'd87;
vramDataLower[12'd1254] = 8'd28;
vramDataLower[12'd1255] = 8'd87;
vramDataLower[12'd1256] = 8'd214;
vramDataLower[12'd1257] = 8'd55;
vramDataLower[12'd1258] = 8'd210;
vramDataLower[12'd1259] = 8'd55;
vramDataLower[12'd1260] = 8'd16;
vramDataLower[12'd1261] = 8'd55;
vramDataLower[12'd1262] = 8'd114;
vramDataLower[12'd1263] = 8'd119;
vramDataLower[12'd1264] = 8'd32;
vramDataLower[12'd1265] = 8'd167;
vramDataLower[12'd1266] = 8'd207;
vramDataLower[12'd1267] = 8'd55;
vramDataLower[12'd1268] = 8'd31;
vramDataLower[12'd1269] = 8'd55;
vramDataLower[12'd1270] = 8'd214;
vramDataLower[12'd1271] = 8'd135;
vramDataLower[12'd1272] = 8'd16;
vramDataLower[12'd1273] = 8'd135;
vramDataLower[12'd1274] = 8'd214;
vramDataLower[12'd1275] = 8'd135;
vramDataLower[12'd1276] = 8'd95;
vramDataLower[12'd1277] = 8'd135;
vramDataLower[12'd1278] = 8'd95;
vramDataLower[12'd1279] = 8'd135;
vramDataLower[12'd1280] = 8'd210;
vramDataLower[12'd1281] = 8'd24;
vramDataLower[12'd1282] = 8'd16;
vramDataLower[12'd1283] = 8'd8;
vramDataLower[12'd1284] = 8'd230;
vramDataLower[12'd1285] = 8'd135;
vramDataLower[12'd1286] = 8'd252;
vramDataLower[12'd1287] = 8'd247;
vramDataLower[12'd1288] = 8'd200;
vramDataLower[12'd1289] = 8'd247;
vramDataLower[12'd1290] = 8'd202;
vramDataLower[12'd1291] = 8'd247;
vramDataLower[12'd1292] = 8'd202;
vramDataLower[12'd1293] = 8'd247;
vramDataLower[12'd1294] = 8'd202;
vramDataLower[12'd1295] = 8'd247;
vramDataLower[12'd1296] = 8'd202;
vramDataLower[12'd1297] = 8'd247;
vramDataLower[12'd1298] = 8'd202;
vramDataLower[12'd1299] = 8'd247;
vramDataLower[12'd1300] = 8'd202;
vramDataLower[12'd1301] = 8'd247;
vramDataLower[12'd1302] = 8'd31;
vramDataLower[12'd1303] = 8'd247;
vramDataLower[12'd1304] = 8'd255;
vramDataLower[12'd1305] = 8'd231;
vramDataLower[12'd1306] = 8'd213;
vramDataLower[12'd1307] = 8'd87;
vramDataLower[12'd1308] = 8'd16;
vramDataLower[12'd1309] = 8'd120;
vramDataLower[12'd1310] = 8'd16;
vramDataLower[12'd1311] = 8'd152;
vramDataLower[12'd1312] = 8'd94;
vramDataLower[12'd1313] = 8'd8;
vramDataLower[12'd1314] = 8'd73;
vramDataLower[12'd1315] = 8'd8;
vramDataLower[12'd1316] = 8'd95;
vramDataLower[12'd1317] = 8'd120;
vramDataLower[12'd1318] = 8'd46;
vramDataLower[12'd1319] = 8'd8;
vramDataLower[12'd1320] = 8'd171;
vramDataLower[12'd1321] = 8'd168;
vramDataLower[12'd1322] = 8'd135;
vramDataLower[12'd1323] = 8'd120;
vramDataLower[12'd1324] = 8'd17;
vramDataLower[12'd1325] = 8'd120;
vramDataLower[12'd1326] = 8'd198;
vramDataLower[12'd1327] = 8'd152;
vramDataLower[12'd1328] = 8'd85;
vramDataLower[12'd1329] = 8'd152;
vramDataLower[12'd1330] = 8'd214;
vramDataLower[12'd1331] = 8'd152;
vramDataLower[12'd1332] = 8'd209;
vramDataLower[12'd1333] = 8'd120;
vramDataLower[12'd1334] = 8'd230;
vramDataLower[12'd1335] = 8'd135;
vramDataLower[12'd1336] = 8'd181;
vramDataLower[12'd1337] = 8'd120;
vramDataLower[12'd1338] = 8'd16;
vramDataLower[12'd1339] = 8'd135;
vramDataLower[12'd1340] = 8'd16;
vramDataLower[12'd1341] = 8'd120;
vramDataLower[12'd1342] = 8'd181;
vramDataLower[12'd1343] = 8'd120;
vramDataLower[12'd1344] = 8'd150;
vramDataLower[12'd1345] = 8'd135;
vramDataLower[12'd1346] = 8'd202;
vramDataLower[12'd1347] = 8'd120;
vramDataLower[12'd1348] = 8'd209;
vramDataLower[12'd1349] = 8'd135;
vramDataLower[12'd1350] = 8'd75;
vramDataLower[12'd1351] = 8'd135;
vramDataLower[12'd1352] = 8'd30;
vramDataLower[12'd1353] = 8'd135;
vramDataLower[12'd1354] = 8'd210;
vramDataLower[12'd1355] = 8'd135;
vramDataLower[12'd1356] = 8'd198;
vramDataLower[12'd1357] = 8'd135;
vramDataLower[12'd1358] = 8'd210;
vramDataLower[12'd1359] = 8'd135;
vramDataLower[12'd1360] = 8'd80;
vramDataLower[12'd1361] = 8'd120;
vramDataLower[12'd1362] = 8'd226;
vramDataLower[12'd1363] = 8'd120;
vramDataLower[12'd1364] = 8'd74;
vramDataLower[12'd1365] = 8'd8;
vramDataLower[12'd1366] = 8'd76;
vramDataLower[12'd1367] = 8'd8;
vramDataLower[12'd1368] = 8'd16;
vramDataLower[12'd1369] = 8'd120;
vramDataLower[12'd1370] = 8'd31;
vramDataLower[12'd1371] = 8'd120;
vramDataLower[12'd1372] = 8'd30;
vramDataLower[12'd1373] = 8'd120;
vramDataLower[12'd1374] = 8'd80;
vramDataLower[12'd1375] = 8'd135;
vramDataLower[12'd1376] = 8'd150;
vramDataLower[12'd1377] = 8'd120;
vramDataLower[12'd1378] = 8'd31;
vramDataLower[12'd1379] = 8'd120;
vramDataLower[12'd1380] = 8'd150;
vramDataLower[12'd1381] = 8'd120;
vramDataLower[12'd1382] = 8'd16;
vramDataLower[12'd1383] = 8'd120;
vramDataLower[12'd1384] = 8'd209;
vramDataLower[12'd1385] = 8'd120;
vramDataLower[12'd1386] = 8'd198;
vramDataLower[12'd1387] = 8'd120;
vramDataLower[12'd1388] = 8'd198;
vramDataLower[12'd1389] = 8'd120;
vramDataLower[12'd1390] = 8'd16;
vramDataLower[12'd1391] = 8'd120;
vramDataLower[12'd1392] = 8'd181;
vramDataLower[12'd1393] = 8'd120;
vramDataLower[12'd1394] = 8'd210;
vramDataLower[12'd1395] = 8'd120;
vramDataLower[12'd1396] = 8'd80;
vramDataLower[12'd1397] = 8'd135;
vramDataLower[12'd1398] = 8'd202;
vramDataLower[12'd1399] = 8'd120;
vramDataLower[12'd1400] = 8'd171;
vramDataLower[12'd1401] = 8'd120;
vramDataLower[12'd1402] = 8'd162;
vramDataLower[12'd1403] = 8'd120;
vramDataLower[12'd1404] = 8'd80;
vramDataLower[12'd1405] = 8'd120;
vramDataLower[12'd1406] = 8'd51;
vramDataLower[12'd1407] = 8'd120;
vramDataLower[12'd1408] = 8'd202;
vramDataLower[12'd1409] = 8'd120;
vramDataLower[12'd1410] = 8'd16;
vramDataLower[12'd1411] = 8'd135;
vramDataLower[12'd1412] = 8'd31;
vramDataLower[12'd1413] = 8'd135;
vramDataLower[12'd1414] = 8'd31;
vramDataLower[12'd1415] = 8'd135;
vramDataLower[12'd1416] = 8'd145;
vramDataLower[12'd1417] = 8'd120;
vramDataLower[12'd1418] = 8'd16;
vramDataLower[12'd1419] = 8'd135;
vramDataLower[12'd1420] = 8'd230;
vramDataLower[12'd1421] = 8'd55;
vramDataLower[12'd1422] = 8'd95;
vramDataLower[12'd1423] = 8'd55;
vramDataLower[12'd1424] = 8'd95;
vramDataLower[12'd1425] = 8'd55;
vramDataLower[12'd1426] = 8'd147;
vramDataLower[12'd1427] = 8'd119;
vramDataLower[12'd1428] = 8'd214;
vramDataLower[12'd1429] = 8'd55;
vramDataLower[12'd1430] = 8'd188;
vramDataLower[12'd1431] = 8'd135;
vramDataLower[12'd1432] = 8'd85;
vramDataLower[12'd1433] = 8'd55;
vramDataLower[12'd1434] = 8'd210;
vramDataLower[12'd1435] = 8'd56;
vramDataLower[12'd1436] = 8'd210;
vramDataLower[12'd1437] = 8'd56;
vramDataLower[12'd1438] = 8'd210;
vramDataLower[12'd1439] = 8'd56;
vramDataLower[12'd1440] = 8'd202;
vramDataLower[12'd1441] = 8'd131;
vramDataLower[12'd1442] = 8'd198;
vramDataLower[12'd1443] = 8'd120;
vramDataLower[12'd1444] = 8'd214;
vramDataLower[12'd1445] = 8'd247;
vramDataLower[12'd1446] = 8'd210;
vramDataLower[12'd1447] = 8'd247;
vramDataLower[12'd1448] = 8'd210;
vramDataLower[12'd1449] = 8'd247;
vramDataLower[12'd1450] = 8'd210;
vramDataLower[12'd1451] = 8'd247;
vramDataLower[12'd1452] = 8'd210;
vramDataLower[12'd1453] = 8'd247;
vramDataLower[12'd1454] = 8'd183;
vramDataLower[12'd1455] = 8'd247;
vramDataLower[12'd1456] = 8'd183;
vramDataLower[12'd1457] = 8'd247;
vramDataLower[12'd1458] = 8'd95;
vramDataLower[12'd1459] = 8'd247;
vramDataLower[12'd1460] = 8'd248;
vramDataLower[12'd1461] = 8'd135;
vramDataLower[12'd1462] = 8'd252;
vramDataLower[12'd1463] = 8'd135;
vramDataLower[12'd1464] = 8'd31;
vramDataLower[12'd1465] = 8'd135;
vramDataLower[12'd1466] = 8'd31;
vramDataLower[12'd1467] = 8'd135;
vramDataLower[12'd1468] = 8'd16;
vramDataLower[12'd1469] = 8'd120;
vramDataLower[12'd1470] = 8'd226;
vramDataLower[12'd1471] = 8'd200;
vramDataLower[12'd1472] = 8'd214;
vramDataLower[12'd1473] = 8'd120;
vramDataLower[12'd1474] = 8'd202;
vramDataLower[12'd1475] = 8'd55;
vramDataLower[12'd1476] = 8'd164;
vramDataLower[12'd1477] = 8'd115;
vramDataLower[12'd1478] = 8'd16;
vramDataLower[12'd1479] = 8'd56;
vramDataLower[12'd1480] = 8'd31;
vramDataLower[12'd1481] = 8'd56;
vramDataLower[12'd1482] = 8'd135;
vramDataLower[12'd1483] = 8'd120;
vramDataLower[12'd1484] = 8'd30;
vramDataLower[12'd1485] = 8'd120;
vramDataLower[12'd1486] = 8'd209;
vramDataLower[12'd1487] = 8'd120;
vramDataLower[12'd1488] = 8'd210;
vramDataLower[12'd1489] = 8'd152;
vramDataLower[12'd1490] = 8'd210;
vramDataLower[12'd1491] = 8'd120;
vramDataLower[12'd1492] = 8'd202;
vramDataLower[12'd1493] = 8'd135;
vramDataLower[12'd1494] = 8'd16;
vramDataLower[12'd1495] = 8'd135;
vramDataLower[12'd1496] = 8'd164;
vramDataLower[12'd1497] = 8'd135;
vramDataLower[12'd1498] = 8'd16;
vramDataLower[12'd1499] = 8'd135;
vramDataLower[12'd1500] = 8'd164;
vramDataLower[12'd1501] = 8'd135;
vramDataLower[12'd1502] = 8'd214;
vramDataLower[12'd1503] = 8'd135;
vramDataLower[12'd1504] = 8'd212;
vramDataLower[12'd1505] = 8'd135;
vramDataLower[12'd1506] = 8'd17;
vramDataLower[12'd1507] = 8'd120;
vramDataLower[12'd1508] = 8'd188;
vramDataLower[12'd1509] = 8'd120;
vramDataLower[12'd1510] = 8'd200;
vramDataLower[12'd1511] = 8'd120;
vramDataLower[12'd1512] = 8'd31;
vramDataLower[12'd1513] = 8'd120;
vramDataLower[12'd1514] = 8'd30;
vramDataLower[12'd1515] = 8'd120;
vramDataLower[12'd1516] = 8'd17;
vramDataLower[12'd1517] = 8'd135;
vramDataLower[12'd1518] = 8'd31;
vramDataLower[12'd1519] = 8'd120;
vramDataLower[12'd1520] = 8'd213;
vramDataLower[12'd1521] = 8'd8;
vramDataLower[12'd1522] = 8'd16;
vramDataLower[12'd1523] = 8'd8;
vramDataLower[12'd1524] = 8'd110;
vramDataLower[12'd1525] = 8'd8;
vramDataLower[12'd1526] = 8'd44;
vramDataLower[12'd1527] = 8'd120;
vramDataLower[12'd1528] = 8'd214;
vramDataLower[12'd1529] = 8'd120;
vramDataLower[12'd1530] = 8'd85;
vramDataLower[12'd1531] = 8'd120;
vramDataLower[12'd1532] = 8'd166;
vramDataLower[12'd1533] = 8'd120;
vramDataLower[12'd1534] = 8'd80;
vramDataLower[12'd1535] = 8'd120;
vramDataLower[12'd1536] = 8'd31;
vramDataLower[12'd1537] = 8'd120;
vramDataLower[12'd1538] = 8'd202;
vramDataLower[12'd1539] = 8'd120;
vramDataLower[12'd1540] = 8'd230;
vramDataLower[12'd1541] = 8'd120;
vramDataLower[12'd1542] = 8'd17;
vramDataLower[12'd1543] = 8'd120;
vramDataLower[12'd1544] = 8'd37;
vramDataLower[12'd1545] = 8'd135;
vramDataLower[12'd1546] = 8'd16;
vramDataLower[12'd1547] = 8'd120;
vramDataLower[12'd1548] = 8'd181;
vramDataLower[12'd1549] = 8'd120;
vramDataLower[12'd1550] = 8'd135;
vramDataLower[12'd1551] = 8'd120;
vramDataLower[12'd1552] = 8'd202;
vramDataLower[12'd1553] = 8'd120;
vramDataLower[12'd1554] = 8'd16;
vramDataLower[12'd1555] = 8'd135;
vramDataLower[12'd1556] = 8'd30;
vramDataLower[12'd1557] = 8'd135;
vramDataLower[12'd1558] = 8'd210;
vramDataLower[12'd1559] = 8'd120;
vramDataLower[12'd1560] = 8'd135;
vramDataLower[12'd1561] = 8'd120;
vramDataLower[12'd1562] = 8'd135;
vramDataLower[12'd1563] = 8'd120;
vramDataLower[12'd1564] = 8'd16;
vramDataLower[12'd1565] = 8'd120;
vramDataLower[12'd1566] = 8'd16;
vramDataLower[12'd1567] = 8'd120;
vramDataLower[12'd1568] = 8'd135;
vramDataLower[12'd1569] = 8'd120;
vramDataLower[12'd1570] = 8'd31;
vramDataLower[12'd1571] = 8'd120;
vramDataLower[12'd1572] = 8'd202;
vramDataLower[12'd1573] = 8'd120;
vramDataLower[12'd1574] = 8'd16;
vramDataLower[12'd1575] = 8'd135;
vramDataLower[12'd1576] = 8'd16;
vramDataLower[12'd1577] = 8'd120;
vramDataLower[12'd1578] = 8'd83;
vramDataLower[12'd1579] = 8'd152;
vramDataLower[12'd1580] = 8'd16;
vramDataLower[12'd1581] = 8'd135;
vramDataLower[12'd1582] = 8'd70;
vramDataLower[12'd1583] = 8'd135;
vramDataLower[12'd1584] = 8'd104;
vramDataLower[12'd1585] = 8'd55;
vramDataLower[12'd1586] = 8'd62;
vramDataLower[12'd1587] = 8'd119;
vramDataLower[12'd1588] = 8'd94;
vramDataLower[12'd1589] = 8'd55;
vramDataLower[12'd1590] = 8'd210;
vramDataLower[12'd1591] = 8'd55;
vramDataLower[12'd1592] = 8'd209;
vramDataLower[12'd1593] = 8'd55;
vramDataLower[12'd1594] = 8'd202;
vramDataLower[12'd1595] = 8'd131;
vramDataLower[12'd1596] = 8'd202;
vramDataLower[12'd1597] = 8'd131;
vramDataLower[12'd1598] = 8'd202;
vramDataLower[12'd1599] = 8'd131;
vramDataLower[12'd1600] = 8'd16;
vramDataLower[12'd1601] = 8'd147;
vramDataLower[12'd1602] = 8'd202;
vramDataLower[12'd1603] = 8'd131;
vramDataLower[12'd1604] = 8'd210;
vramDataLower[12'd1605] = 8'd55;
vramDataLower[12'd1606] = 8'd210;
vramDataLower[12'd1607] = 8'd55;
vramDataLower[12'd1608] = 8'd183;
vramDataLower[12'd1609] = 8'd55;
vramDataLower[12'd1610] = 8'd183;
vramDataLower[12'd1611] = 8'd55;
vramDataLower[12'd1612] = 8'd252;
vramDataLower[12'd1613] = 8'd247;
vramDataLower[12'd1614] = 8'd202;
vramDataLower[12'd1615] = 8'd247;
vramDataLower[12'd1616] = 8'd202;
vramDataLower[12'd1617] = 8'd247;
vramDataLower[12'd1618] = 8'd202;
vramDataLower[12'd1619] = 8'd247;
vramDataLower[12'd1620] = 8'd202;
vramDataLower[12'd1621] = 8'd247;
vramDataLower[12'd1622] = 8'd202;
vramDataLower[12'd1623] = 8'd247;
vramDataLower[12'd1624] = 8'd248;
vramDataLower[12'd1625] = 8'd247;
vramDataLower[12'd1626] = 8'd214;
vramDataLower[12'd1627] = 8'd135;
vramDataLower[12'd1628] = 8'd80;
vramDataLower[12'd1629] = 8'd120;
vramDataLower[12'd1630] = 8'd239;
vramDataLower[12'd1631] = 8'd152;
vramDataLower[12'd1632] = 8'd145;
vramDataLower[12'd1633] = 8'd55;
vramDataLower[12'd1634] = 8'd209;
vramDataLower[12'd1635] = 8'd55;
vramDataLower[12'd1636] = 8'd202;
vramDataLower[12'd1637] = 8'd55;
vramDataLower[12'd1638] = 8'd198;
vramDataLower[12'd1639] = 8'd8;
vramDataLower[12'd1640] = 8'd213;
vramDataLower[12'd1641] = 8'd56;
vramDataLower[12'd1642] = 8'd164;
vramDataLower[12'd1643] = 8'd55;
vramDataLower[12'd1644] = 8'd16;
vramDataLower[12'd1645] = 8'd120;
vramDataLower[12'd1646] = 8'd16;
vramDataLower[12'd1647] = 8'd120;
vramDataLower[12'd1648] = 8'd164;
vramDataLower[12'd1649] = 8'd135;
vramDataLower[12'd1650] = 8'd30;
vramDataLower[12'd1651] = 8'd135;
vramDataLower[12'd1652] = 8'd164;
vramDataLower[12'd1653] = 8'd135;
vramDataLower[12'd1654] = 8'd16;
vramDataLower[12'd1655] = 8'd135;
vramDataLower[12'd1656] = 8'd124;
vramDataLower[12'd1657] = 8'd135;
vramDataLower[12'd1658] = 8'd17;
vramDataLower[12'd1659] = 8'd135;
vramDataLower[12'd1660] = 8'd124;
vramDataLower[12'd1661] = 8'd135;
vramDataLower[12'd1662] = 8'd102;
vramDataLower[12'd1663] = 8'd135;
vramDataLower[12'd1664] = 8'd124;
vramDataLower[12'd1665] = 8'd135;
vramDataLower[12'd1666] = 8'd252;
vramDataLower[12'd1667] = 8'd135;
vramDataLower[12'd1668] = 8'd16;
vramDataLower[12'd1669] = 8'd120;
vramDataLower[12'd1670] = 8'd230;
vramDataLower[12'd1671] = 8'd120;
vramDataLower[12'd1672] = 8'd109;
vramDataLower[12'd1673] = 8'd120;
vramDataLower[12'd1674] = 8'd195;
vramDataLower[12'd1675] = 8'd152;
vramDataLower[12'd1676] = 8'd198;
vramDataLower[12'd1677] = 8'd120;
vramDataLower[12'd1678] = 8'd250;
vramDataLower[12'd1679] = 8'd8;
vramDataLower[12'd1680] = 8'd200;
vramDataLower[12'd1681] = 8'd8;
vramDataLower[12'd1682] = 8'd73;
vramDataLower[12'd1683] = 8'd8;
vramDataLower[12'd1684] = 8'd61;
vramDataLower[12'd1685] = 8'd152;
vramDataLower[12'd1686] = 8'd17;
vramDataLower[12'd1687] = 8'd152;
vramDataLower[12'd1688] = 8'd55;
vramDataLower[12'd1689] = 8'd120;
vramDataLower[12'd1690] = 8'd159;
vramDataLower[12'd1691] = 8'd120;
vramDataLower[12'd1692] = 8'd228;
vramDataLower[12'd1693] = 8'd120;
vramDataLower[12'd1694] = 8'd30;
vramDataLower[12'd1695] = 8'd120;
vramDataLower[12'd1696] = 8'd135;
vramDataLower[12'd1697] = 8'd120;
vramDataLower[12'd1698] = 8'd210;
vramDataLower[12'd1699] = 8'd120;
vramDataLower[12'd1700] = 8'd51;
vramDataLower[12'd1701] = 8'd120;
vramDataLower[12'd1702] = 8'd253;
vramDataLower[12'd1703] = 8'd135;
vramDataLower[12'd1704] = 8'd95;
vramDataLower[12'd1705] = 8'd135;
vramDataLower[12'd1706] = 8'd50;
vramDataLower[12'd1707] = 8'd135;
vramDataLower[12'd1708] = 8'd209;
vramDataLower[12'd1709] = 8'd135;
vramDataLower[12'd1710] = 8'd83;
vramDataLower[12'd1711] = 8'd120;
vramDataLower[12'd1712] = 8'd159;
vramDataLower[12'd1713] = 8'd120;
vramDataLower[12'd1714] = 8'd202;
vramDataLower[12'd1715] = 8'd120;
vramDataLower[12'd1716] = 8'd202;
vramDataLower[12'd1717] = 8'd120;
vramDataLower[12'd1718] = 8'd148;
vramDataLower[12'd1719] = 8'd120;
vramDataLower[12'd1720] = 8'd30;
vramDataLower[12'd1721] = 8'd120;
vramDataLower[12'd1722] = 8'd50;
vramDataLower[12'd1723] = 8'd120;
vramDataLower[12'd1724] = 8'd210;
vramDataLower[12'd1725] = 8'd120;
vramDataLower[12'd1726] = 8'd202;
vramDataLower[12'd1727] = 8'd120;
vramDataLower[12'd1728] = 8'd172;
vramDataLower[12'd1729] = 8'd120;
vramDataLower[12'd1730] = 8'd166;
vramDataLower[12'd1731] = 8'd120;
vramDataLower[12'd1732] = 8'd17;
vramDataLower[12'd1733] = 8'd120;
vramDataLower[12'd1734] = 8'd150;
vramDataLower[12'd1735] = 8'd120;
vramDataLower[12'd1736] = 8'd16;
vramDataLower[12'd1737] = 8'd120;
vramDataLower[12'd1738] = 8'd210;
vramDataLower[12'd1739] = 8'd120;
vramDataLower[12'd1740] = 8'd210;
vramDataLower[12'd1741] = 8'd135;
vramDataLower[12'd1742] = 8'd16;
vramDataLower[12'd1743] = 8'd135;
vramDataLower[12'd1744] = 8'd95;
vramDataLower[12'd1745] = 8'd55;
vramDataLower[12'd1746] = 8'd95;
vramDataLower[12'd1747] = 8'd55;
vramDataLower[12'd1748] = 8'd200;
vramDataLower[12'd1749] = 8'd55;
vramDataLower[12'd1750] = 8'd164;
vramDataLower[12'd1751] = 8'd55;
vramDataLower[12'd1752] = 8'd80;
vramDataLower[12'd1753] = 8'd115;
vramDataLower[12'd1754] = 8'd145;
vramDataLower[12'd1755] = 8'd131;
vramDataLower[12'd1756] = 8'd202;
vramDataLower[12'd1757] = 8'd131;
vramDataLower[12'd1758] = 8'd202;
vramDataLower[12'd1759] = 8'd131;
vramDataLower[12'd1760] = 8'd202;
vramDataLower[12'd1761] = 8'd147;
vramDataLower[12'd1762] = 8'd202;
vramDataLower[12'd1763] = 8'd147;
vramDataLower[12'd1764] = 8'd202;
vramDataLower[12'd1765] = 8'd147;
vramDataLower[12'd1766] = 8'd202;
vramDataLower[12'd1767] = 8'd115;
vramDataLower[12'd1768] = 8'd210;
vramDataLower[12'd1769] = 8'd55;
vramDataLower[12'd1770] = 8'd210;
vramDataLower[12'd1771] = 8'd55;
vramDataLower[12'd1772] = 8'd210;
vramDataLower[12'd1773] = 8'd55;
vramDataLower[12'd1774] = 8'd210;
vramDataLower[12'd1775] = 8'd55;
vramDataLower[12'd1776] = 8'd210;
vramDataLower[12'd1777] = 8'd55;
vramDataLower[12'd1778] = 8'd210;
vramDataLower[12'd1779] = 8'd55;
vramDataLower[12'd1780] = 8'd181;
vramDataLower[12'd1781] = 8'd55;
vramDataLower[12'd1782] = 8'd16;
vramDataLower[12'd1783] = 8'd55;
vramDataLower[12'd1784] = 8'd30;
vramDataLower[12'd1785] = 8'd135;
vramDataLower[12'd1786] = 8'd31;
vramDataLower[12'd1787] = 8'd135;
vramDataLower[12'd1788] = 8'd226;
vramDataLower[12'd1789] = 8'd120;
vramDataLower[12'd1790] = 8'd17;
vramDataLower[12'd1791] = 8'd8;
vramDataLower[12'd1792] = 8'd16;
vramDataLower[12'd1793] = 8'd55;
vramDataLower[12'd1794] = 8'd202;
vramDataLower[12'd1795] = 8'd55;
vramDataLower[12'd1796] = 8'd210;
vramDataLower[12'd1797] = 8'd55;
vramDataLower[12'd1798] = 8'd16;
vramDataLower[12'd1799] = 8'd135;
vramDataLower[12'd1800] = 8'd31;
vramDataLower[12'd1801] = 8'd247;
vramDataLower[12'd1802] = 8'd80;
vramDataLower[12'd1803] = 8'd55;
vramDataLower[12'd1804] = 8'd17;
vramDataLower[12'd1805] = 8'd135;
vramDataLower[12'd1806] = 8'd181;
vramDataLower[12'd1807] = 8'd135;
vramDataLower[12'd1808] = 8'd181;
vramDataLower[12'd1809] = 8'd135;
vramDataLower[12'd1810] = 8'd188;
vramDataLower[12'd1811] = 8'd135;
vramDataLower[12'd1812] = 8'd34;
vramDataLower[12'd1813] = 8'd55;
vramDataLower[12'd1814] = 8'd58;
vramDataLower[12'd1815] = 8'd247;
vramDataLower[12'd1816] = 8'd239;
vramDataLower[12'd1817] = 8'd135;
vramDataLower[12'd1818] = 8'd76;
vramDataLower[12'd1819] = 8'd247;
vramDataLower[12'd1820] = 8'd170;
vramDataLower[12'd1821] = 8'd135;
vramDataLower[12'd1822] = 8'd89;
vramDataLower[12'd1823] = 8'd247;
vramDataLower[12'd1824] = 8'd96;
vramDataLower[12'd1825] = 8'd247;
vramDataLower[12'd1826] = 8'd218;
vramDataLower[12'd1827] = 8'd135;
vramDataLower[12'd1828] = 8'd96;
vramDataLower[12'd1829] = 8'd135;
vramDataLower[12'd1830] = 8'd104;
vramDataLower[12'd1831] = 8'd135;
vramDataLower[12'd1832] = 8'd190;
vramDataLower[12'd1833] = 8'd135;
vramDataLower[12'd1834] = 8'd200;
vramDataLower[12'd1835] = 8'd135;
vramDataLower[12'd1836] = 8'd16;
vramDataLower[12'd1837] = 8'd120;
vramDataLower[12'd1838] = 8'd16;
vramDataLower[12'd1839] = 8'd120;
vramDataLower[12'd1840] = 8'd16;
vramDataLower[12'd1841] = 8'd152;
vramDataLower[12'd1842] = 8'd127;
vramDataLower[12'd1843] = 8'd120;
vramDataLower[12'd1844] = 8'd248;
vramDataLower[12'd1845] = 8'd120;
vramDataLower[12'd1846] = 8'd30;
vramDataLower[12'd1847] = 8'd120;
vramDataLower[12'd1848] = 8'd30;
vramDataLower[12'd1849] = 8'd120;
vramDataLower[12'd1850] = 8'd202;
vramDataLower[12'd1851] = 8'd120;
vramDataLower[12'd1852] = 8'd202;
vramDataLower[12'd1853] = 8'd120;
vramDataLower[12'd1854] = 8'd30;
vramDataLower[12'd1855] = 8'd135;
vramDataLower[12'd1856] = 8'd155;
vramDataLower[12'd1857] = 8'd135;
vramDataLower[12'd1858] = 8'd31;
vramDataLower[12'd1859] = 8'd135;
vramDataLower[12'd1860] = 8'd202;
vramDataLower[12'd1861] = 8'd135;
vramDataLower[12'd1862] = 8'd51;
vramDataLower[12'd1863] = 8'd135;
vramDataLower[12'd1864] = 8'd16;
vramDataLower[12'd1865] = 8'd135;
vramDataLower[12'd1866] = 8'd30;
vramDataLower[12'd1867] = 8'd135;
vramDataLower[12'd1868] = 8'd31;
vramDataLower[12'd1869] = 8'd135;
vramDataLower[12'd1870] = 8'd202;
vramDataLower[12'd1871] = 8'd135;
vramDataLower[12'd1872] = 8'd17;
vramDataLower[12'd1873] = 8'd120;
vramDataLower[12'd1874] = 8'd210;
vramDataLower[12'd1875] = 8'd120;
vramDataLower[12'd1876] = 8'd135;
vramDataLower[12'd1877] = 8'd120;
vramDataLower[12'd1878] = 8'd208;
vramDataLower[12'd1879] = 8'd120;
vramDataLower[12'd1880] = 8'd207;
vramDataLower[12'd1881] = 8'd120;
vramDataLower[12'd1882] = 8'd164;
vramDataLower[12'd1883] = 8'd120;
vramDataLower[12'd1884] = 8'd31;
vramDataLower[12'd1885] = 8'd120;
vramDataLower[12'd1886] = 8'd31;
vramDataLower[12'd1887] = 8'd120;
vramDataLower[12'd1888] = 8'd16;
vramDataLower[12'd1889] = 8'd120;
vramDataLower[12'd1890] = 8'd95;
vramDataLower[12'd1891] = 8'd120;
vramDataLower[12'd1892] = 8'd95;
vramDataLower[12'd1893] = 8'd120;
vramDataLower[12'd1894] = 8'd208;
vramDataLower[12'd1895] = 8'd120;
vramDataLower[12'd1896] = 8'd30;
vramDataLower[12'd1897] = 8'd120;
vramDataLower[12'd1898] = 8'd135;
vramDataLower[12'd1899] = 8'd152;
vramDataLower[12'd1900] = 8'd214;
vramDataLower[12'd1901] = 8'd120;
vramDataLower[12'd1902] = 8'd210;
vramDataLower[12'd1903] = 8'd120;
vramDataLower[12'd1904] = 8'd16;
vramDataLower[12'd1905] = 8'd120;
vramDataLower[12'd1906] = 8'd16;
vramDataLower[12'd1907] = 8'd135;
vramDataLower[12'd1908] = 8'd17;
vramDataLower[12'd1909] = 8'd247;
vramDataLower[12'd1910] = 8'd214;
vramDataLower[12'd1911] = 8'd55;
vramDataLower[12'd1912] = 8'd164;
vramDataLower[12'd1913] = 8'd131;
vramDataLower[12'd1914] = 8'd202;
vramDataLower[12'd1915] = 8'd131;
vramDataLower[12'd1916] = 8'd210;
vramDataLower[12'd1917] = 8'd131;
vramDataLower[12'd1918] = 8'd202;
vramDataLower[12'd1919] = 8'd131;
vramDataLower[12'd1920] = 8'd202;
vramDataLower[12'd1921] = 8'd147;
vramDataLower[12'd1922] = 8'd202;
vramDataLower[12'd1923] = 8'd147;
vramDataLower[12'd1924] = 8'd202;
vramDataLower[12'd1925] = 8'd147;
vramDataLower[12'd1926] = 8'd202;
vramDataLower[12'd1927] = 8'd147;
vramDataLower[12'd1928] = 8'd202;
vramDataLower[12'd1929] = 8'd147;
vramDataLower[12'd1930] = 8'd202;
vramDataLower[12'd1931] = 8'd147;
vramDataLower[12'd1932] = 8'd202;
vramDataLower[12'd1933] = 8'd147;
vramDataLower[12'd1934] = 8'd202;
vramDataLower[12'd1935] = 8'd147;
vramDataLower[12'd1936] = 8'd202;
vramDataLower[12'd1937] = 8'd147;
vramDataLower[12'd1938] = 8'd202;
vramDataLower[12'd1939] = 8'd147;
vramDataLower[12'd1940] = 8'd210;
vramDataLower[12'd1941] = 8'd135;
vramDataLower[12'd1942] = 8'd164;
vramDataLower[12'd1943] = 8'd120;
vramDataLower[12'd1944] = 8'd16;
vramDataLower[12'd1945] = 8'd135;
vramDataLower[12'd1946] = 8'd209;
vramDataLower[12'd1947] = 8'd135;
vramDataLower[12'd1948] = 8'd16;
vramDataLower[12'd1949] = 8'd120;
vramDataLower[12'd1950] = 8'd200;
vramDataLower[12'd1951] = 8'd8;
vramDataLower[12'd1952] = 8'd30;
vramDataLower[12'd1953] = 8'd8;
vramDataLower[12'd1954] = 8'd202;
vramDataLower[12'd1955] = 8'd56;
vramDataLower[12'd1956] = 8'd202;
vramDataLower[12'd1957] = 8'd115;
vramDataLower[12'd1958] = 8'd210;
vramDataLower[12'd1959] = 8'd55;
vramDataLower[12'd1960] = 8'd210;
vramDataLower[12'd1961] = 8'd55;
vramDataLower[12'd1962] = 8'd198;
vramDataLower[12'd1963] = 8'd135;
vramDataLower[12'd1964] = 8'd214;
vramDataLower[12'd1965] = 8'd135;
vramDataLower[12'd1966] = 8'd145;
vramDataLower[12'd1967] = 8'd135;
vramDataLower[12'd1968] = 8'd135;
vramDataLower[12'd1969] = 8'd135;
vramDataLower[12'd1970] = 8'd104;
vramDataLower[12'd1971] = 8'd135;
vramDataLower[12'd1972] = 8'd7;
vramDataLower[12'd1973] = 8'd247;
vramDataLower[12'd1974] = 8'd28;
vramDataLower[12'd1975] = 8'd135;
vramDataLower[12'd1976] = 8'd164;
vramDataLower[12'd1977] = 8'd247;
vramDataLower[12'd1978] = 8'd109;
vramDataLower[12'd1979] = 8'd247;
vramDataLower[12'd1980] = 8'd9;
vramDataLower[12'd1981] = 8'd247;
vramDataLower[12'd1982] = 8'd39;
vramDataLower[12'd1983] = 8'd247;
vramDataLower[12'd1984] = 8'd24;
vramDataLower[12'd1985] = 8'd103;
vramDataLower[12'd1986] = 8'd16;
vramDataLower[12'd1987] = 8'd247;
vramDataLower[12'd1988] = 8'd17;
vramDataLower[12'd1989] = 8'd247;
vramDataLower[12'd1990] = 8'd17;
vramDataLower[12'd1991] = 8'd247;
vramDataLower[12'd1992] = 8'd95;
vramDataLower[12'd1993] = 8'd247;
vramDataLower[12'd1994] = 8'd39;
vramDataLower[12'd1995] = 8'd135;
vramDataLower[12'd1996] = 8'd16;
vramDataLower[12'd1997] = 8'd120;
vramDataLower[12'd1998] = 8'd80;
vramDataLower[12'd1999] = 8'd120;
vramDataLower[12'd2000] = 8'd94;
vramDataLower[12'd2001] = 8'd152;
vramDataLower[12'd2002] = 8'd214;
vramDataLower[12'd2003] = 8'd8;
vramDataLower[12'd2004] = 8'd31;
vramDataLower[12'd2005] = 8'd8;
vramDataLower[12'd2006] = 8'd202;
vramDataLower[12'd2007] = 8'd8;
vramDataLower[12'd2008] = 8'd95;
vramDataLower[12'd2009] = 8'd56;
vramDataLower[12'd2010] = 8'd214;
vramDataLower[12'd2011] = 8'd152;
vramDataLower[12'd2012] = 8'd95;
vramDataLower[12'd2013] = 8'd56;
vramDataLower[12'd2014] = 8'd95;
vramDataLower[12'd2015] = 8'd56;
vramDataLower[12'd2016] = 8'd95;
vramDataLower[12'd2017] = 8'd56;
vramDataLower[12'd2018] = 8'd126;
vramDataLower[12'd2019] = 8'd120;
vramDataLower[12'd2020] = 8'd200;
vramDataLower[12'd2021] = 8'd120;
vramDataLower[12'd2022] = 8'd30;
vramDataLower[12'd2023] = 8'd120;
vramDataLower[12'd2024] = 8'd83;
vramDataLower[12'd2025] = 8'd120;
vramDataLower[12'd2026] = 8'd239;
vramDataLower[12'd2027] = 8'd135;
vramDataLower[12'd2028] = 8'd167;
vramDataLower[12'd2029] = 8'd135;
vramDataLower[12'd2030] = 8'd166;
vramDataLower[12'd2031] = 8'd135;
vramDataLower[12'd2032] = 8'd226;
vramDataLower[12'd2033] = 8'd135;
vramDataLower[12'd2034] = 8'd240;
vramDataLower[12'd2035] = 8'd120;
vramDataLower[12'd2036] = 8'd17;
vramDataLower[12'd2037] = 8'd120;
vramDataLower[12'd2038] = 8'd80;
vramDataLower[12'd2039] = 8'd120;
vramDataLower[12'd2040] = 8'd181;
vramDataLower[12'd2041] = 8'd120;
vramDataLower[12'd2042] = 8'd37;
vramDataLower[12'd2043] = 8'd120;
vramDataLower[12'd2044] = 8'd16;
vramDataLower[12'd2045] = 8'd120;
vramDataLower[12'd2046] = 8'd31;
vramDataLower[12'd2047] = 8'd120;
vramDataLower[12'd2048] = 8'd83;
vramDataLower[12'd2049] = 8'd120;
vramDataLower[12'd2050] = 8'd210;
vramDataLower[12'd2051] = 8'd120;
vramDataLower[12'd2052] = 8'd17;
vramDataLower[12'd2053] = 8'd120;
vramDataLower[12'd2054] = 8'd202;
vramDataLower[12'd2055] = 8'd120;
vramDataLower[12'd2056] = 8'd31;
vramDataLower[12'd2057] = 8'd120;
vramDataLower[12'd2058] = 8'd70;
vramDataLower[12'd2059] = 8'd120;
vramDataLower[12'd2060] = 8'd208;
vramDataLower[12'd2061] = 8'd120;
vramDataLower[12'd2062] = 8'd210;
vramDataLower[12'd2063] = 8'd120;
vramDataLower[12'd2064] = 8'd223;
vramDataLower[12'd2065] = 8'd135;
vramDataLower[12'd2066] = 8'd214;
vramDataLower[12'd2067] = 8'd55;
vramDataLower[12'd2068] = 8'd80;
vramDataLower[12'd2069] = 8'd120;
vramDataLower[12'd2070] = 8'd202;
vramDataLower[12'd2071] = 8'd56;
vramDataLower[12'd2072] = 8'd202;
vramDataLower[12'd2073] = 8'd56;
vramDataLower[12'd2074] = 8'd202;
vramDataLower[12'd2075] = 8'd56;
vramDataLower[12'd2076] = 8'd202;
vramDataLower[12'd2077] = 8'd56;
vramDataLower[12'd2078] = 8'd202;
vramDataLower[12'd2079] = 8'd56;
vramDataLower[12'd2080] = 8'd202;
vramDataLower[12'd2081] = 8'd24;
vramDataLower[12'd2082] = 8'd202;
vramDataLower[12'd2083] = 8'd24;
vramDataLower[12'd2084] = 8'd202;
vramDataLower[12'd2085] = 8'd24;
vramDataLower[12'd2086] = 8'd202;
vramDataLower[12'd2087] = 8'd24;
vramDataLower[12'd2088] = 8'd202;
vramDataLower[12'd2089] = 8'd24;
vramDataLower[12'd2090] = 8'd210;
vramDataLower[12'd2091] = 8'd8;
vramDataLower[12'd2092] = 8'd210;
vramDataLower[12'd2093] = 8'd8;
vramDataLower[12'd2094] = 8'd16;
vramDataLower[12'd2095] = 8'd8;
vramDataLower[12'd2096] = 8'd202;
vramDataLower[12'd2097] = 8'd56;
vramDataLower[12'd2098] = 8'd202;
vramDataLower[12'd2099] = 8'd56;
vramDataLower[12'd2100] = 8'd80;
vramDataLower[12'd2101] = 8'd152;
vramDataLower[12'd2102] = 8'd202;
vramDataLower[12'd2103] = 8'd152;
vramDataLower[12'd2104] = 8'd202;
vramDataLower[12'd2105] = 8'd152;
vramDataLower[12'd2106] = 8'd51;
vramDataLower[12'd2107] = 8'd120;
vramDataLower[12'd2108] = 8'd210;
vramDataLower[12'd2109] = 8'd135;
vramDataLower[12'd2110] = 8'd208;
vramDataLower[12'd2111] = 8'd135;
vramDataLower[12'd2112] = 8'd202;
vramDataLower[12'd2113] = 8'd135;
vramDataLower[12'd2114] = 8'd220;
vramDataLower[12'd2115] = 8'd120;
vramDataLower[12'd2116] = 8'd210;
vramDataLower[12'd2117] = 8'd120;
vramDataLower[12'd2118] = 8'd210;
vramDataLower[12'd2119] = 8'd120;
vramDataLower[12'd2120] = 8'd31;
vramDataLower[12'd2121] = 8'd135;
vramDataLower[12'd2122] = 8'd31;
vramDataLower[12'd2123] = 8'd135;
vramDataLower[12'd2124] = 8'd220;
vramDataLower[12'd2125] = 8'd120;
vramDataLower[12'd2126] = 8'd253;
vramDataLower[12'd2127] = 8'd135;
vramDataLower[12'd2128] = 8'd205;
vramDataLower[12'd2129] = 8'd135;
vramDataLower[12'd2130] = 8'd95;
vramDataLower[12'd2131] = 8'd247;
vramDataLower[12'd2132] = 8'd89;
vramDataLower[12'd2133] = 8'd247;
vramDataLower[12'd2134] = 8'd202;
vramDataLower[12'd2135] = 8'd247;
vramDataLower[12'd2136] = 8'd19;
vramDataLower[12'd2137] = 8'd247;
vramDataLower[12'd2138] = 8'd89;
vramDataLower[12'd2139] = 8'd247;
vramDataLower[12'd2140] = 8'd93;
vramDataLower[12'd2141] = 8'd247;
vramDataLower[12'd2142] = 8'd245;
vramDataLower[12'd2143] = 8'd247;
vramDataLower[12'd2144] = 8'd200;
vramDataLower[12'd2145] = 8'd247;
vramDataLower[12'd2146] = 8'd129;
vramDataLower[12'd2147] = 8'd247;
vramDataLower[12'd2148] = 8'd30;
vramDataLower[12'd2149] = 8'd247;
vramDataLower[12'd2150] = 8'd86;
vramDataLower[12'd2151] = 8'd247;
vramDataLower[12'd2152] = 8'd33;
vramDataLower[12'd2153] = 8'd87;
vramDataLower[12'd2154] = 8'd31;
vramDataLower[12'd2155] = 8'd135;
vramDataLower[12'd2156] = 8'd171;
vramDataLower[12'd2157] = 8'd120;
vramDataLower[12'd2158] = 8'd95;
vramDataLower[12'd2159] = 8'd8;
vramDataLower[12'd2160] = 8'd214;
vramDataLower[12'd2161] = 8'd8;
vramDataLower[12'd2162] = 8'd16;
vramDataLower[12'd2163] = 8'd8;
vramDataLower[12'd2164] = 8'd80;
vramDataLower[12'd2165] = 8'd135;
vramDataLower[12'd2166] = 8'd202;
vramDataLower[12'd2167] = 8'd55;
vramDataLower[12'd2168] = 8'd202;
vramDataLower[12'd2169] = 8'd55;
vramDataLower[12'd2170] = 8'd31;
vramDataLower[12'd2171] = 8'd115;
vramDataLower[12'd2172] = 8'd16;
vramDataLower[12'd2173] = 8'd120;
vramDataLower[12'd2174] = 8'd31;
vramDataLower[12'd2175] = 8'd8;
vramDataLower[12'd2176] = 8'd198;
vramDataLower[12'd2177] = 8'd120;
vramDataLower[12'd2178] = 8'd16;
vramDataLower[12'd2179] = 8'd55;
vramDataLower[12'd2180] = 8'd209;
vramDataLower[12'd2181] = 8'd55;
vramDataLower[12'd2182] = 8'd183;
vramDataLower[12'd2183] = 8'd120;
vramDataLower[12'd2184] = 8'd230;
vramDataLower[12'd2185] = 8'd152;
vramDataLower[12'd2186] = 8'd200;
vramDataLower[12'd2187] = 8'd120;
vramDataLower[12'd2188] = 8'd83;
vramDataLower[12'd2189] = 8'd135;
vramDataLower[12'd2190] = 8'd16;
vramDataLower[12'd2191] = 8'd135;
vramDataLower[12'd2192] = 8'd50;
vramDataLower[12'd2193] = 8'd135;
vramDataLower[12'd2194] = 8'd80;
vramDataLower[12'd2195] = 8'd135;
vramDataLower[12'd2196] = 8'd17;
vramDataLower[12'd2197] = 8'd120;
vramDataLower[12'd2198] = 8'd198;
vramDataLower[12'd2199] = 8'd120;
vramDataLower[12'd2200] = 8'd210;
vramDataLower[12'd2201] = 8'd120;
vramDataLower[12'd2202] = 8'd80;
vramDataLower[12'd2203] = 8'd120;
vramDataLower[12'd2204] = 8'd51;
vramDataLower[12'd2205] = 8'd120;
vramDataLower[12'd2206] = 8'd156;
vramDataLower[12'd2207] = 8'd120;
vramDataLower[12'd2208] = 8'd51;
vramDataLower[12'd2209] = 8'd120;
vramDataLower[12'd2210] = 8'd17;
vramDataLower[12'd2211] = 8'd120;
vramDataLower[12'd2212] = 8'd214;
vramDataLower[12'd2213] = 8'd120;
vramDataLower[12'd2214] = 8'd17;
vramDataLower[12'd2215] = 8'd120;
vramDataLower[12'd2216] = 8'd202;
vramDataLower[12'd2217] = 8'd120;
vramDataLower[12'd2218] = 8'd171;
vramDataLower[12'd2219] = 8'd120;
vramDataLower[12'd2220] = 8'd214;
vramDataLower[12'd2221] = 8'd120;
vramDataLower[12'd2222] = 8'd226;
vramDataLower[12'd2223] = 8'd135;
vramDataLower[12'd2224] = 8'd226;
vramDataLower[12'd2225] = 8'd247;
vramDataLower[12'd2226] = 8'd198;
vramDataLower[12'd2227] = 8'd55;
vramDataLower[12'd2228] = 8'd16;
vramDataLower[12'd2229] = 8'd147;
vramDataLower[12'd2230] = 8'd202;
vramDataLower[12'd2231] = 8'd19;
vramDataLower[12'd2232] = 8'd202;
vramDataLower[12'd2233] = 8'd19;
vramDataLower[12'd2234] = 8'd202;
vramDataLower[12'd2235] = 8'd19;
vramDataLower[12'd2236] = 8'd202;
vramDataLower[12'd2237] = 8'd19;
vramDataLower[12'd2238] = 8'd202;
vramDataLower[12'd2239] = 8'd19;
vramDataLower[12'd2240] = 8'd210;
vramDataLower[12'd2241] = 8'd115;
vramDataLower[12'd2242] = 8'd202;
vramDataLower[12'd2243] = 8'd131;
vramDataLower[12'd2244] = 8'd202;
vramDataLower[12'd2245] = 8'd131;
vramDataLower[12'd2246] = 8'd210;
vramDataLower[12'd2247] = 8'd56;
vramDataLower[12'd2248] = 8'd164;
vramDataLower[12'd2249] = 8'd24;
vramDataLower[12'd2250] = 8'd202;
vramDataLower[12'd2251] = 8'd24;
vramDataLower[12'd2252] = 8'd80;
vramDataLower[12'd2253] = 8'd8;
vramDataLower[12'd2254] = 8'd95;
vramDataLower[12'd2255] = 8'd8;
vramDataLower[12'd2256] = 8'd202;
vramDataLower[12'd2257] = 8'd152;
vramDataLower[12'd2258] = 8'd202;
vramDataLower[12'd2259] = 8'd152;
vramDataLower[12'd2260] = 8'd202;
vramDataLower[12'd2261] = 8'd152;
vramDataLower[12'd2262] = 8'd135;
vramDataLower[12'd2263] = 8'd152;
vramDataLower[12'd2264] = 8'd202;
vramDataLower[12'd2265] = 8'd152;
vramDataLower[12'd2266] = 8'd109;
vramDataLower[12'd2267] = 8'd152;
vramDataLower[12'd2268] = 8'd166;
vramDataLower[12'd2269] = 8'd120;
vramDataLower[12'd2270] = 8'd16;
vramDataLower[12'd2271] = 8'd135;
vramDataLower[12'd2272] = 8'd135;
vramDataLower[12'd2273] = 8'd135;
vramDataLower[12'd2274] = 8'd16;
vramDataLower[12'd2275] = 8'd135;
vramDataLower[12'd2276] = 8'd31;
vramDataLower[12'd2277] = 8'd55;
vramDataLower[12'd2278] = 8'd80;
vramDataLower[12'd2279] = 8'd55;
vramDataLower[12'd2280] = 8'd183;
vramDataLower[12'd2281] = 8'd247;
vramDataLower[12'd2282] = 8'd51;
vramDataLower[12'd2283] = 8'd247;
vramDataLower[12'd2284] = 8'd226;
vramDataLower[12'd2285] = 8'd247;
vramDataLower[12'd2286] = 8'd70;
vramDataLower[12'd2287] = 8'd247;
vramDataLower[12'd2288] = 8'd52;
vramDataLower[12'd2289] = 8'd247;
vramDataLower[12'd2290] = 8'd167;
vramDataLower[12'd2291] = 8'd247;
vramDataLower[12'd2292] = 8'd107;
vramDataLower[12'd2293] = 8'd247;
vramDataLower[12'd2294] = 8'd119;
vramDataLower[12'd2295] = 8'd247;
vramDataLower[12'd2296] = 8'd190;
vramDataLower[12'd2297] = 8'd247;
vramDataLower[12'd2298] = 8'd16;
vramDataLower[12'd2299] = 8'd247;
vramDataLower[12'd2300] = 8'd16;
vramDataLower[12'd2301] = 8'd247;
vramDataLower[12'd2302] = 8'd30;
vramDataLower[12'd2303] = 8'd247;
vramDataLower[12'd2304] = 8'd156;
vramDataLower[12'd2305] = 8'd247;
vramDataLower[12'd2306] = 8'd202;
vramDataLower[12'd2307] = 8'd247;
vramDataLower[12'd2308] = 8'd75;
vramDataLower[12'd2309] = 8'd247;
vramDataLower[12'd2310] = 8'd24;
vramDataLower[12'd2311] = 8'd87;
vramDataLower[12'd2312] = 8'd218;
vramDataLower[12'd2313] = 8'd247;
vramDataLower[12'd2314] = 8'd226;
vramDataLower[12'd2315] = 8'd120;
vramDataLower[12'd2316] = 8'd210;
vramDataLower[12'd2317] = 8'd8;
vramDataLower[12'd2318] = 8'd37;
vramDataLower[12'd2319] = 8'd128;
vramDataLower[12'd2320] = 8'd164;
vramDataLower[12'd2321] = 8'd8;
vramDataLower[12'd2322] = 8'd221;
vramDataLower[12'd2323] = 8'd135;
vramDataLower[12'd2324] = 8'd209;
vramDataLower[12'd2325] = 8'd183;
vramDataLower[12'd2326] = 8'd16;
vramDataLower[12'd2327] = 8'd183;
vramDataLower[12'd2328] = 8'd17;
vramDataLower[12'd2329] = 8'd183;
vramDataLower[12'd2330] = 8'd16;
vramDataLower[12'd2331] = 8'd183;
vramDataLower[12'd2332] = 8'd16;
vramDataLower[12'd2333] = 8'd8;
vramDataLower[12'd2334] = 8'd16;
vramDataLower[12'd2335] = 8'd8;
vramDataLower[12'd2336] = 8'd80;
vramDataLower[12'd2337] = 8'd135;
vramDataLower[12'd2338] = 8'd80;
vramDataLower[12'd2339] = 8'd183;
vramDataLower[12'd2340] = 8'd16;
vramDataLower[12'd2341] = 8'd183;
vramDataLower[12'd2342] = 8'd31;
vramDataLower[12'd2343] = 8'd247;
vramDataLower[12'd2344] = 8'd200;
vramDataLower[12'd2345] = 8'd55;
vramDataLower[12'd2346] = 8'd16;
vramDataLower[12'd2347] = 8'd120;
vramDataLower[12'd2348] = 8'd17;
vramDataLower[12'd2349] = 8'd120;
vramDataLower[12'd2350] = 8'd16;
vramDataLower[12'd2351] = 8'd135;
vramDataLower[12'd2352] = 8'd164;
vramDataLower[12'd2353] = 8'd135;
vramDataLower[12'd2354] = 8'd83;
vramDataLower[12'd2355] = 8'd120;
vramDataLower[12'd2356] = 8'd209;
vramDataLower[12'd2357] = 8'd120;
vramDataLower[12'd2358] = 8'd37;
vramDataLower[12'd2359] = 8'd135;
vramDataLower[12'd2360] = 8'd202;
vramDataLower[12'd2361] = 8'd135;
vramDataLower[12'd2362] = 8'd31;
vramDataLower[12'd2363] = 8'd120;
vramDataLower[12'd2364] = 8'd197;
vramDataLower[12'd2365] = 8'd120;
vramDataLower[12'd2366] = 8'd9;
vramDataLower[12'd2367] = 8'd120;
vramDataLower[12'd2368] = 8'd31;
vramDataLower[12'd2369] = 8'd135;
vramDataLower[12'd2370] = 8'd31;
vramDataLower[12'd2371] = 8'd135;
vramDataLower[12'd2372] = 8'd61;
vramDataLower[12'd2373] = 8'd135;
vramDataLower[12'd2374] = 8'd200;
vramDataLower[12'd2375] = 8'd135;
vramDataLower[12'd2376] = 8'd202;
vramDataLower[12'd2377] = 8'd135;
vramDataLower[12'd2378] = 8'd202;
vramDataLower[12'd2379] = 8'd135;
vramDataLower[12'd2380] = 8'd253;
vramDataLower[12'd2381] = 8'd135;
vramDataLower[12'd2382] = 8'd75;
vramDataLower[12'd2383] = 8'd119;
vramDataLower[12'd2384] = 8'd16;
vramDataLower[12'd2385] = 8'd87;
vramDataLower[12'd2386] = 8'd198;
vramDataLower[12'd2387] = 8'd55;
vramDataLower[12'd2388] = 8'd210;
vramDataLower[12'd2389] = 8'd147;
vramDataLower[12'd2390] = 8'd16;
vramDataLower[12'd2391] = 8'd147;
vramDataLower[12'd2392] = 8'd210;
vramDataLower[12'd2393] = 8'd147;
vramDataLower[12'd2394] = 8'd210;
vramDataLower[12'd2395] = 8'd147;
vramDataLower[12'd2396] = 8'd210;
vramDataLower[12'd2397] = 8'd147;
vramDataLower[12'd2398] = 8'd210;
vramDataLower[12'd2399] = 8'd147;
vramDataLower[12'd2400] = 8'd210;
vramDataLower[12'd2401] = 8'd147;
vramDataLower[12'd2402] = 8'd210;
vramDataLower[12'd2403] = 8'd147;
vramDataLower[12'd2404] = 8'd210;
vramDataLower[12'd2405] = 8'd147;
vramDataLower[12'd2406] = 8'd202;
vramDataLower[12'd2407] = 8'd131;
vramDataLower[12'd2408] = 8'd16;
vramDataLower[12'd2409] = 8'd56;
vramDataLower[12'd2410] = 8'd145;
vramDataLower[12'd2411] = 8'd24;
vramDataLower[12'd2412] = 8'd202;
vramDataLower[12'd2413] = 8'd8;
vramDataLower[12'd2414] = 8'd31;
vramDataLower[12'd2415] = 8'd8;
vramDataLower[12'd2416] = 8'd16;
vramDataLower[12'd2417] = 8'd8;
vramDataLower[12'd2418] = 8'd214;
vramDataLower[12'd2419] = 8'd152;
vramDataLower[12'd2420] = 8'd181;
vramDataLower[12'd2421] = 8'd152;
vramDataLower[12'd2422] = 8'd85;
vramDataLower[12'd2423] = 8'd152;
vramDataLower[12'd2424] = 8'd210;
vramDataLower[12'd2425] = 8'd152;
vramDataLower[12'd2426] = 8'd214;
vramDataLower[12'd2427] = 8'd120;
vramDataLower[12'd2428] = 8'd80;
vramDataLower[12'd2429] = 8'd135;
vramDataLower[12'd2430] = 8'd202;
vramDataLower[12'd2431] = 8'd135;
vramDataLower[12'd2432] = 8'd31;
vramDataLower[12'd2433] = 8'd55;
vramDataLower[12'd2434] = 8'd202;
vramDataLower[12'd2435] = 8'd55;
vramDataLower[12'd2436] = 8'd248;
vramDataLower[12'd2437] = 8'd55;
vramDataLower[12'd2438] = 8'd37;
vramDataLower[12'd2439] = 8'd247;
vramDataLower[12'd2440] = 8'd230;
vramDataLower[12'd2441] = 8'd247;
vramDataLower[12'd2442] = 8'd241;
vramDataLower[12'd2443] = 8'd247;
vramDataLower[12'd2444] = 8'd210;
vramDataLower[12'd2445] = 8'd247;
vramDataLower[12'd2446] = 8'd240;
vramDataLower[12'd2447] = 8'd247;
vramDataLower[12'd2448] = 8'd171;
vramDataLower[12'd2449] = 8'd247;
vramDataLower[12'd2450] = 8'd31;
vramDataLower[12'd2451] = 8'd247;
vramDataLower[12'd2452] = 8'd86;
vramDataLower[12'd2453] = 8'd247;
vramDataLower[12'd2454] = 8'd106;
vramDataLower[12'd2455] = 8'd247;
vramDataLower[12'd2456] = 8'd181;
vramDataLower[12'd2457] = 8'd247;
vramDataLower[12'd2458] = 8'd7;
vramDataLower[12'd2459] = 8'd247;
vramDataLower[12'd2460] = 8'd239;
vramDataLower[12'd2461] = 8'd247;
vramDataLower[12'd2462] = 8'd252;
vramDataLower[12'd2463] = 8'd247;
vramDataLower[12'd2464] = 8'd198;
vramDataLower[12'd2465] = 8'd87;
vramDataLower[12'd2466] = 8'd31;
vramDataLower[12'd2467] = 8'd135;
vramDataLower[12'd2468] = 8'd240;
vramDataLower[12'd2469] = 8'd247;
vramDataLower[12'd2470] = 8'd218;
vramDataLower[12'd2471] = 8'd247;
vramDataLower[12'd2472] = 8'd188;
vramDataLower[12'd2473] = 8'd247;
vramDataLower[12'd2474] = 8'd202;
vramDataLower[12'd2475] = 8'd135;
vramDataLower[12'd2476] = 8'd200;
vramDataLower[12'd2477] = 8'd8;
vramDataLower[12'd2478] = 8'd16;
vramDataLower[12'd2479] = 8'd128;
vramDataLower[12'd2480] = 8'd17;
vramDataLower[12'd2481] = 8'd128;
vramDataLower[12'd2482] = 8'd200;
vramDataLower[12'd2483] = 8'd120;
vramDataLower[12'd2484] = 8'd202;
vramDataLower[12'd2485] = 8'd183;
vramDataLower[12'd2486] = 8'd164;
vramDataLower[12'd2487] = 8'd183;
vramDataLower[12'd2488] = 8'd209;
vramDataLower[12'd2489] = 8'd183;
vramDataLower[12'd2490] = 8'd181;
vramDataLower[12'd2491] = 8'd183;
vramDataLower[12'd2492] = 8'd223;
vramDataLower[12'd2493] = 8'd135;
vramDataLower[12'd2494] = 8'd70;
vramDataLower[12'd2495] = 8'd135;
vramDataLower[12'd2496] = 8'd37;
vramDataLower[12'd2497] = 8'd247;
vramDataLower[12'd2498] = 8'd30;
vramDataLower[12'd2499] = 8'd183;
vramDataLower[12'd2500] = 8'd210;
vramDataLower[12'd2501] = 8'd183;
vramDataLower[12'd2502] = 8'd16;
vramDataLower[12'd2503] = 8'd183;
vramDataLower[12'd2504] = 8'd220;
vramDataLower[12'd2505] = 8'd135;
vramDataLower[12'd2506] = 8'd76;
vramDataLower[12'd2507] = 8'd152;
vramDataLower[12'd2508] = 8'd67;
vramDataLower[12'd2509] = 8'd135;
vramDataLower[12'd2510] = 8'd17;
vramDataLower[12'd2511] = 8'd135;
vramDataLower[12'd2512] = 8'd171;
vramDataLower[12'd2513] = 8'd120;
vramDataLower[12'd2514] = 8'd202;
vramDataLower[12'd2515] = 8'd120;
vramDataLower[12'd2516] = 8'd117;
vramDataLower[12'd2517] = 8'd120;
vramDataLower[12'd2518] = 8'd37;
vramDataLower[12'd2519] = 8'd120;
vramDataLower[12'd2520] = 8'd30;
vramDataLower[12'd2521] = 8'd135;
vramDataLower[12'd2522] = 8'd240;
vramDataLower[12'd2523] = 8'd120;
vramDataLower[12'd2524] = 8'd156;
vramDataLower[12'd2525] = 8'd135;
vramDataLower[12'd2526] = 8'd240;
vramDataLower[12'd2527] = 8'd135;
vramDataLower[12'd2528] = 8'd240;
vramDataLower[12'd2529] = 8'd135;
vramDataLower[12'd2530] = 8'd30;
vramDataLower[12'd2531] = 8'd135;
vramDataLower[12'd2532] = 8'd17;
vramDataLower[12'd2533] = 8'd135;
vramDataLower[12'd2534] = 8'd46;
vramDataLower[12'd2535] = 8'd135;
vramDataLower[12'd2536] = 8'd126;
vramDataLower[12'd2537] = 8'd135;
vramDataLower[12'd2538] = 8'd135;
vramDataLower[12'd2539] = 8'd55;
vramDataLower[12'd2540] = 8'd16;
vramDataLower[12'd2541] = 8'd55;
vramDataLower[12'd2542] = 8'd71;
vramDataLower[12'd2543] = 8'd119;
vramDataLower[12'd2544] = 8'd117;
vramDataLower[12'd2545] = 8'd247;
vramDataLower[12'd2546] = 8'd16;
vramDataLower[12'd2547] = 8'd247;
vramDataLower[12'd2548] = 8'd16;
vramDataLower[12'd2549] = 8'd115;
vramDataLower[12'd2550] = 8'd145;
vramDataLower[12'd2551] = 8'd179;
vramDataLower[12'd2552] = 8'd145;
vramDataLower[12'd2553] = 8'd179;
vramDataLower[12'd2554] = 8'd145;
vramDataLower[12'd2555] = 8'd179;
vramDataLower[12'd2556] = 8'd145;
vramDataLower[12'd2557] = 8'd179;
vramDataLower[12'd2558] = 8'd16;
vramDataLower[12'd2559] = 8'd179;
vramDataLower[12'd2560] = 8'd210;
vramDataLower[12'd2561] = 8'd147;
vramDataLower[12'd2562] = 8'd181;
vramDataLower[12'd2563] = 8'd147;
vramDataLower[12'd2564] = 8'd202;
vramDataLower[12'd2565] = 8'd147;
vramDataLower[12'd2566] = 8'd164;
vramDataLower[12'd2567] = 8'd147;
vramDataLower[12'd2568] = 8'd202;
vramDataLower[12'd2569] = 8'd131;
vramDataLower[12'd2570] = 8'd202;
vramDataLower[12'd2571] = 8'd131;
vramDataLower[12'd2572] = 8'd145;
vramDataLower[12'd2573] = 8'd24;
vramDataLower[12'd2574] = 8'd214;
vramDataLower[12'd2575] = 8'd152;
vramDataLower[12'd2576] = 8'd70;
vramDataLower[12'd2577] = 8'd135;
vramDataLower[12'd2578] = 8'd200;
vramDataLower[12'd2579] = 8'd135;
vramDataLower[12'd2580] = 8'd16;
vramDataLower[12'd2581] = 8'd120;
vramDataLower[12'd2582] = 8'd210;
vramDataLower[12'd2583] = 8'd120;
vramDataLower[12'd2584] = 8'd210;
vramDataLower[12'd2585] = 8'd120;
vramDataLower[12'd2586] = 8'd16;
vramDataLower[12'd2587] = 8'd135;
vramDataLower[12'd2588] = 8'd164;
vramDataLower[12'd2589] = 8'd55;
vramDataLower[12'd2590] = 8'd30;
vramDataLower[12'd2591] = 8'd55;
vramDataLower[12'd2592] = 8'd214;
vramDataLower[12'd2593] = 8'd247;
vramDataLower[12'd2594] = 8'd9;
vramDataLower[12'd2595] = 8'd247;
vramDataLower[12'd2596] = 8'd107;
vramDataLower[12'd2597] = 8'd247;
vramDataLower[12'd2598] = 8'd241;
vramDataLower[12'd2599] = 8'd247;
vramDataLower[12'd2600] = 8'd31;
vramDataLower[12'd2601] = 8'd247;
vramDataLower[12'd2602] = 8'd157;
vramDataLower[12'd2603] = 8'd247;
vramDataLower[12'd2604] = 8'd83;
vramDataLower[12'd2605] = 8'd247;
vramDataLower[12'd2606] = 8'd83;
vramDataLower[12'd2607] = 8'd247;
vramDataLower[12'd2608] = 8'd37;
vramDataLower[12'd2609] = 8'd247;
vramDataLower[12'd2610] = 8'd109;
vramDataLower[12'd2611] = 8'd247;
vramDataLower[12'd2612] = 8'd108;
vramDataLower[12'd2613] = 8'd247;
vramDataLower[12'd2614] = 8'd252;
vramDataLower[12'd2615] = 8'd247;
vramDataLower[12'd2616] = 8'd159;
vramDataLower[12'd2617] = 8'd247;
vramDataLower[12'd2618] = 8'd86;
vramDataLower[12'd2619] = 8'd247;
vramDataLower[12'd2620] = 8'd95;
vramDataLower[12'd2621] = 8'd135;
vramDataLower[12'd2622] = 8'd52;
vramDataLower[12'd2623] = 8'd135;
vramDataLower[12'd2624] = 8'd52;
vramDataLower[12'd2625] = 8'd135;
vramDataLower[12'd2626] = 8'd16;
vramDataLower[12'd2627] = 8'd135;
vramDataLower[12'd2628] = 8'd127;
vramDataLower[12'd2629] = 8'd135;
vramDataLower[12'd2630] = 8'd28;
vramDataLower[12'd2631] = 8'd135;
vramDataLower[12'd2632] = 8'd183;
vramDataLower[12'd2633] = 8'd87;
vramDataLower[12'd2634] = 8'd16;
vramDataLower[12'd2635] = 8'd87;
vramDataLower[12'd2636] = 8'd46;
vramDataLower[12'd2637] = 8'd135;
vramDataLower[12'd2638] = 8'd200;
vramDataLower[12'd2639] = 8'd135;
vramDataLower[12'd2640] = 8'd183;
vramDataLower[12'd2641] = 8'd120;
vramDataLower[12'd2642] = 8'd166;
vramDataLower[12'd2643] = 8'd8;
vramDataLower[12'd2644] = 8'd202;
vramDataLower[12'd2645] = 8'd56;
vramDataLower[12'd2646] = 8'd223;
vramDataLower[12'd2647] = 8'd120;
vramDataLower[12'd2648] = 8'd145;
vramDataLower[12'd2649] = 8'd183;
vramDataLower[12'd2650] = 8'd145;
vramDataLower[12'd2651] = 8'd183;
vramDataLower[12'd2652] = 8'd210;
vramDataLower[12'd2653] = 8'd55;
vramDataLower[12'd2654] = 8'd210;
vramDataLower[12'd2655] = 8'd55;
vramDataLower[12'd2656] = 8'd210;
vramDataLower[12'd2657] = 8'd55;
vramDataLower[12'd2658] = 8'd202;
vramDataLower[12'd2659] = 8'd115;
vramDataLower[12'd2660] = 8'd80;
vramDataLower[12'd2661] = 8'd56;
vramDataLower[12'd2662] = 8'd95;
vramDataLower[12'd2663] = 8'd120;
vramDataLower[12'd2664] = 8'd214;
vramDataLower[12'd2665] = 8'd120;
vramDataLower[12'd2666] = 8'd107;
vramDataLower[12'd2667] = 8'd135;
vramDataLower[12'd2668] = 8'd164;
vramDataLower[12'd2669] = 8'd135;
vramDataLower[12'd2670] = 8'd67;
vramDataLower[12'd2671] = 8'd135;
vramDataLower[12'd2672] = 8'd18;
vramDataLower[12'd2673] = 8'd135;
vramDataLower[12'd2674] = 8'd210;
vramDataLower[12'd2675] = 8'd135;
vramDataLower[12'd2676] = 8'd210;
vramDataLower[12'd2677] = 8'd120;
vramDataLower[12'd2678] = 8'd210;
vramDataLower[12'd2679] = 8'd120;
vramDataLower[12'd2680] = 8'd30;
vramDataLower[12'd2681] = 8'd120;
vramDataLower[12'd2682] = 8'd90;
vramDataLower[12'd2683] = 8'd120;
vramDataLower[12'd2684] = 8'd101;
vramDataLower[12'd2685] = 8'd120;
vramDataLower[12'd2686] = 8'd240;
vramDataLower[12'd2687] = 8'd135;
vramDataLower[12'd2688] = 8'd240;
vramDataLower[12'd2689] = 8'd135;
vramDataLower[12'd2690] = 8'd240;
vramDataLower[12'd2691] = 8'd135;
vramDataLower[12'd2692] = 8'd28;
vramDataLower[12'd2693] = 8'd135;
vramDataLower[12'd2694] = 8'd226;
vramDataLower[12'd2695] = 8'd135;
vramDataLower[12'd2696] = 8'd51;
vramDataLower[12'd2697] = 8'd55;
vramDataLower[12'd2698] = 8'd31;
vramDataLower[12'd2699] = 8'd55;
vramDataLower[12'd2700] = 8'd92;
vramDataLower[12'd2701] = 8'd55;
vramDataLower[12'd2702] = 8'd95;
vramDataLower[12'd2703] = 8'd247;
vramDataLower[12'd2704] = 8'd192;
vramDataLower[12'd2705] = 8'd119;
vramDataLower[12'd2706] = 8'd30;
vramDataLower[12'd2707] = 8'd247;
vramDataLower[12'd2708] = 8'd222;
vramDataLower[12'd2709] = 8'd135;
vramDataLower[12'd2710] = 8'd202;
vramDataLower[12'd2711] = 8'd56;
vramDataLower[12'd2712] = 8'd223;
vramDataLower[12'd2713] = 8'd56;
vramDataLower[12'd2714] = 8'd220;
vramDataLower[12'd2715] = 8'd131;
vramDataLower[12'd2716] = 8'd220;
vramDataLower[12'd2717] = 8'd131;
vramDataLower[12'd2718] = 8'd220;
vramDataLower[12'd2719] = 8'd131;
vramDataLower[12'd2720] = 8'd202;
vramDataLower[12'd2721] = 8'd147;
vramDataLower[12'd2722] = 8'd202;
vramDataLower[12'd2723] = 8'd147;
vramDataLower[12'd2724] = 8'd181;
vramDataLower[12'd2725] = 8'd147;
vramDataLower[12'd2726] = 8'd210;
vramDataLower[12'd2727] = 8'd147;
vramDataLower[12'd2728] = 8'd210;
vramDataLower[12'd2729] = 8'd147;
vramDataLower[12'd2730] = 8'd202;
vramDataLower[12'd2731] = 8'd131;
vramDataLower[12'd2732] = 8'd210;
vramDataLower[12'd2733] = 8'd56;
vramDataLower[12'd2734] = 8'd70;
vramDataLower[12'd2735] = 8'd55;
vramDataLower[12'd2736] = 8'd183;
vramDataLower[12'd2737] = 8'd247;
vramDataLower[12'd2738] = 8'd95;
vramDataLower[12'd2739] = 8'd247;
vramDataLower[12'd2740] = 8'd200;
vramDataLower[12'd2741] = 8'd135;
vramDataLower[12'd2742] = 8'd202;
vramDataLower[12'd2743] = 8'd135;
vramDataLower[12'd2744] = 8'd210;
vramDataLower[12'd2745] = 8'd135;
vramDataLower[12'd2746] = 8'd210;
vramDataLower[12'd2747] = 8'd55;
vramDataLower[12'd2748] = 8'd230;
vramDataLower[12'd2749] = 8'd55;
vramDataLower[12'd2750] = 8'd95;
vramDataLower[12'd2751] = 8'd135;
vramDataLower[12'd2752] = 8'd210;
vramDataLower[12'd2753] = 8'd55;
vramDataLower[12'd2754] = 8'd28;
vramDataLower[12'd2755] = 8'd55;
vramDataLower[12'd2756] = 8'd228;
vramDataLower[12'd2757] = 8'd55;
vramDataLower[12'd2758] = 8'd253;
vramDataLower[12'd2759] = 8'd247;
vramDataLower[12'd2760] = 8'd162;
vramDataLower[12'd2761] = 8'd247;
vramDataLower[12'd2762] = 8'd197;
vramDataLower[12'd2763] = 8'd247;
vramDataLower[12'd2764] = 8'd202;
vramDataLower[12'd2765] = 8'd247;
vramDataLower[12'd2766] = 8'd239;
vramDataLower[12'd2767] = 8'd247;
vramDataLower[12'd2768] = 8'd202;
vramDataLower[12'd2769] = 8'd247;
vramDataLower[12'd2770] = 8'd252;
vramDataLower[12'd2771] = 8'd247;
vramDataLower[12'd2772] = 8'd253;
vramDataLower[12'd2773] = 8'd247;
vramDataLower[12'd2774] = 8'd102;
vramDataLower[12'd2775] = 8'd135;
vramDataLower[12'd2776] = 8'd253;
vramDataLower[12'd2777] = 8'd247;
vramDataLower[12'd2778] = 8'd212;
vramDataLower[12'd2779] = 8'd135;
vramDataLower[12'd2780] = 8'd30;
vramDataLower[12'd2781] = 8'd135;
vramDataLower[12'd2782] = 8'd107;
vramDataLower[12'd2783] = 8'd135;
vramDataLower[12'd2784] = 8'd252;
vramDataLower[12'd2785] = 8'd135;
vramDataLower[12'd2786] = 8'd16;
vramDataLower[12'd2787] = 8'd135;
vramDataLower[12'd2788] = 8'd115;
vramDataLower[12'd2789] = 8'd135;
vramDataLower[12'd2790] = 8'd26;
vramDataLower[12'd2791] = 8'd135;
vramDataLower[12'd2792] = 8'd16;
vramDataLower[12'd2793] = 8'd135;
vramDataLower[12'd2794] = 8'd34;
vramDataLower[12'd2795] = 8'd135;
vramDataLower[12'd2796] = 8'd50;
vramDataLower[12'd2797] = 8'd135;
vramDataLower[12'd2798] = 8'd228;
vramDataLower[12'd2799] = 8'd135;
vramDataLower[12'd2800] = 8'd118;
vramDataLower[12'd2801] = 8'd135;
vramDataLower[12'd2802] = 8'd162;
vramDataLower[12'd2803] = 8'd135;
vramDataLower[12'd2804] = 8'd200;
vramDataLower[12'd2805] = 8'd135;
vramDataLower[12'd2806] = 8'd208;
vramDataLower[12'd2807] = 8'd135;
vramDataLower[12'd2808] = 8'd220;
vramDataLower[12'd2809] = 8'd120;
vramDataLower[12'd2810] = 8'd223;
vramDataLower[12'd2811] = 8'd135;
vramDataLower[12'd2812] = 8'd223;
vramDataLower[12'd2813] = 8'd135;
vramDataLower[12'd2814] = 8'd17;
vramDataLower[12'd2815] = 8'd120;
vramDataLower[12'd2816] = 8'd223;
vramDataLower[12'd2817] = 8'd135;
vramDataLower[12'd2818] = 8'd202;
vramDataLower[12'd2819] = 8'd135;
vramDataLower[12'd2820] = 8'd83;
vramDataLower[12'd2821] = 8'd135;
vramDataLower[12'd2822] = 8'd17;
vramDataLower[12'd2823] = 8'd135;
vramDataLower[12'd2824] = 8'd135;
vramDataLower[12'd2825] = 8'd135;
vramDataLower[12'd2826] = 8'd228;
vramDataLower[12'd2827] = 8'd135;
vramDataLower[12'd2828] = 8'd101;
vramDataLower[12'd2829] = 8'd135;
vramDataLower[12'd2830] = 8'd149;
vramDataLower[12'd2831] = 8'd135;
vramDataLower[12'd2832] = 8'd52;
vramDataLower[12'd2833] = 8'd135;
vramDataLower[12'd2834] = 8'd9;
vramDataLower[12'd2835] = 8'd135;
vramDataLower[12'd2836] = 8'd16;
vramDataLower[12'd2837] = 8'd135;
vramDataLower[12'd2838] = 8'd209;
vramDataLower[12'd2839] = 8'd135;
vramDataLower[12'd2840] = 8'd70;
vramDataLower[12'd2841] = 8'd135;
vramDataLower[12'd2842] = 8'd209;
vramDataLower[12'd2843] = 8'd135;
vramDataLower[12'd2844] = 8'd83;
vramDataLower[12'd2845] = 8'd135;
vramDataLower[12'd2846] = 8'd95;
vramDataLower[12'd2847] = 8'd135;
vramDataLower[12'd2848] = 8'd37;
vramDataLower[12'd2849] = 8'd135;
vramDataLower[12'd2850] = 8'd31;
vramDataLower[12'd2851] = 8'd135;
vramDataLower[12'd2852] = 8'd240;
vramDataLower[12'd2853] = 8'd135;
vramDataLower[12'd2854] = 8'd76;
vramDataLower[12'd2855] = 8'd87;
vramDataLower[12'd2856] = 8'd95;
vramDataLower[12'd2857] = 8'd135;
vramDataLower[12'd2858] = 8'd240;
vramDataLower[12'd2859] = 8'd55;
vramDataLower[12'd2860] = 8'd28;
vramDataLower[12'd2861] = 8'd55;
vramDataLower[12'd2862] = 8'd212;
vramDataLower[12'd2863] = 8'd247;
vramDataLower[12'd2864] = 8'd135;
vramDataLower[12'd2865] = 8'd247;
vramDataLower[12'd2866] = 8'd18;
vramDataLower[12'd2867] = 8'd247;
vramDataLower[12'd2868] = 8'd16;
vramDataLower[12'd2869] = 8'd120;
vramDataLower[12'd2870] = 8'd122;
vramDataLower[12'd2871] = 8'd152;
vramDataLower[12'd2872] = 8'd198;
vramDataLower[12'd2873] = 8'd24;
vramDataLower[12'd2874] = 8'd209;
vramDataLower[12'd2875] = 8'd24;
vramDataLower[12'd2876] = 8'd210;
vramDataLower[12'd2877] = 8'd24;
vramDataLower[12'd2878] = 8'd210;
vramDataLower[12'd2879] = 8'd16;
vramDataLower[12'd2880] = 8'd202;
vramDataLower[12'd2881] = 8'd147;
vramDataLower[12'd2882] = 8'd202;
vramDataLower[12'd2883] = 8'd147;
vramDataLower[12'd2884] = 8'd210;
vramDataLower[12'd2885] = 8'd147;
vramDataLower[12'd2886] = 8'd202;
vramDataLower[12'd2887] = 8'd147;
vramDataLower[12'd2888] = 8'd83;
vramDataLower[12'd2889] = 8'd147;
vramDataLower[12'd2890] = 8'd210;
vramDataLower[12'd2891] = 8'd147;
vramDataLower[12'd2892] = 8'd70;
vramDataLower[12'd2893] = 8'd55;
vramDataLower[12'd2894] = 8'd145;
vramDataLower[12'd2895] = 8'd247;
vramDataLower[12'd2896] = 8'd145;
vramDataLower[12'd2897] = 8'd247;
vramDataLower[12'd2898] = 8'd16;
vramDataLower[12'd2899] = 8'd247;
vramDataLower[12'd2900] = 8'd197;
vramDataLower[12'd2901] = 8'd135;
vramDataLower[12'd2902] = 8'd253;
vramDataLower[12'd2903] = 8'd120;
vramDataLower[12'd2904] = 8'd200;
vramDataLower[12'd2905] = 8'd152;
vramDataLower[12'd2906] = 8'd202;
vramDataLower[12'd2907] = 8'd120;
vramDataLower[12'd2908] = 8'd214;
vramDataLower[12'd2909] = 8'd135;
vramDataLower[12'd2910] = 8'd135;
vramDataLower[12'd2911] = 8'd135;
vramDataLower[12'd2912] = 8'd209;
vramDataLower[12'd2913] = 8'd135;
vramDataLower[12'd2914] = 8'd210;
vramDataLower[12'd2915] = 8'd135;
vramDataLower[12'd2916] = 8'd135;
vramDataLower[12'd2917] = 8'd135;
vramDataLower[12'd2918] = 8'd51;
vramDataLower[12'd2919] = 8'd87;
vramDataLower[12'd2920] = 8'd96;
vramDataLower[12'd2921] = 8'd247;
vramDataLower[12'd2922] = 8'd208;
vramDataLower[12'd2923] = 8'd247;
vramDataLower[12'd2924] = 8'd9;
vramDataLower[12'd2925] = 8'd247;
vramDataLower[12'd2926] = 8'd9;
vramDataLower[12'd2927] = 8'd247;
vramDataLower[12'd2928] = 8'd46;
vramDataLower[12'd2929] = 8'd135;
vramDataLower[12'd2930] = 8'd191;
vramDataLower[12'd2931] = 8'd135;
vramDataLower[12'd2932] = 8'd59;
vramDataLower[12'd2933] = 8'd247;
vramDataLower[12'd2934] = 8'd95;
vramDataLower[12'd2935] = 8'd135;
vramDataLower[12'd2936] = 8'd126;
vramDataLower[12'd2937] = 8'd135;
vramDataLower[12'd2938] = 8'd250;
vramDataLower[12'd2939] = 8'd247;
vramDataLower[12'd2940] = 8'd164;
vramDataLower[12'd2941] = 8'd135;
vramDataLower[12'd2942] = 8'd200;
vramDataLower[12'd2943] = 8'd135;
vramDataLower[12'd2944] = 8'd30;
vramDataLower[12'd2945] = 8'd135;
vramDataLower[12'd2946] = 8'd122;
vramDataLower[12'd2947] = 8'd135;
vramDataLower[12'd2948] = 8'd92;
vramDataLower[12'd2949] = 8'd135;
vramDataLower[12'd2950] = 8'd89;
vramDataLower[12'd2951] = 8'd135;
vramDataLower[12'd2952] = 8'd253;
vramDataLower[12'd2953] = 8'd135;
vramDataLower[12'd2954] = 8'd210;
vramDataLower[12'd2955] = 8'd135;
vramDataLower[12'd2956] = 8'd17;
vramDataLower[12'd2957] = 8'd120;
vramDataLower[12'd2958] = 8'd88;
vramDataLower[12'd2959] = 8'd135;
vramDataLower[12'd2960] = 8'd210;
vramDataLower[12'd2961] = 8'd135;
vramDataLower[12'd2962] = 8'd171;
vramDataLower[12'd2963] = 8'd135;
vramDataLower[12'd2964] = 8'd210;
vramDataLower[12'd2965] = 8'd135;
vramDataLower[12'd2966] = 8'd97;
vramDataLower[12'd2967] = 8'd135;
vramDataLower[12'd2968] = 8'd83;
vramDataLower[12'd2969] = 8'd120;
vramDataLower[12'd2970] = 8'd83;
vramDataLower[12'd2971] = 8'd120;
vramDataLower[12'd2972] = 8'd228;
vramDataLower[12'd2973] = 8'd120;
vramDataLower[12'd2974] = 8'd208;
vramDataLower[12'd2975] = 8'd120;
vramDataLower[12'd2976] = 8'd200;
vramDataLower[12'd2977] = 8'd120;
vramDataLower[12'd2978] = 8'd80;
vramDataLower[12'd2979] = 8'd120;
vramDataLower[12'd2980] = 8'd228;
vramDataLower[12'd2981] = 8'd120;
vramDataLower[12'd2982] = 8'd248;
vramDataLower[12'd2983] = 8'd120;
vramDataLower[12'd2984] = 8'd226;
vramDataLower[12'd2985] = 8'd120;
vramDataLower[12'd2986] = 8'd164;
vramDataLower[12'd2987] = 8'd120;
vramDataLower[12'd2988] = 8'd171;
vramDataLower[12'd2989] = 8'd120;
vramDataLower[12'd2990] = 8'd198;
vramDataLower[12'd2991] = 8'd120;
vramDataLower[12'd2992] = 8'd31;
vramDataLower[12'd2993] = 8'd120;
vramDataLower[12'd2994] = 8'd31;
vramDataLower[12'd2995] = 8'd120;
vramDataLower[12'd2996] = 8'd240;
vramDataLower[12'd2997] = 8'd135;
vramDataLower[12'd2998] = 8'd210;
vramDataLower[12'd2999] = 8'd135;
vramDataLower[12'd3000] = 8'd16;
vramDataLower[12'd3001] = 8'd135;
vramDataLower[12'd3002] = 8'd30;
vramDataLower[12'd3003] = 8'd135;
vramDataLower[12'd3004] = 8'd239;
vramDataLower[12'd3005] = 8'd135;
vramDataLower[12'd3006] = 8'd102;
vramDataLower[12'd3007] = 8'd135;
vramDataLower[12'd3008] = 8'd95;
vramDataLower[12'd3009] = 8'd135;
vramDataLower[12'd3010] = 8'd42;
vramDataLower[12'd3011] = 8'd135;
vramDataLower[12'd3012] = 8'd76;
vramDataLower[12'd3013] = 8'd135;
vramDataLower[12'd3014] = 8'd247;
vramDataLower[12'd3015] = 8'd135;
vramDataLower[12'd3016] = 8'd31;
vramDataLower[12'd3017] = 8'd135;
vramDataLower[12'd3018] = 8'd126;
vramDataLower[12'd3019] = 8'd55;
vramDataLower[12'd3020] = 8'd31;
vramDataLower[12'd3021] = 8'd135;
vramDataLower[12'd3022] = 8'd95;
vramDataLower[12'd3023] = 8'd55;
vramDataLower[12'd3024] = 8'd37;
vramDataLower[12'd3025] = 8'd247;
vramDataLower[12'd3026] = 8'd16;
vramDataLower[12'd3027] = 8'd247;
vramDataLower[12'd3028] = 8'd16;
vramDataLower[12'd3029] = 8'd120;
vramDataLower[12'd3030] = 8'd210;
vramDataLower[12'd3031] = 8'd56;
vramDataLower[12'd3032] = 8'd210;
vramDataLower[12'd3033] = 8'd56;
vramDataLower[12'd3034] = 8'd202;
vramDataLower[12'd3035] = 8'd24;
vramDataLower[12'd3036] = 8'd148;
vramDataLower[12'd3037] = 8'd129;
vramDataLower[12'd3038] = 8'd164;
vramDataLower[12'd3039] = 8'd129;
vramDataLower[12'd3040] = 8'd16;
vramDataLower[12'd3041] = 8'd19;
vramDataLower[12'd3042] = 8'd148;
vramDataLower[12'd3043] = 8'd147;
vramDataLower[12'd3044] = 8'd83;
vramDataLower[12'd3045] = 8'd147;
vramDataLower[12'd3046] = 8'd202;
vramDataLower[12'd3047] = 8'd147;
vramDataLower[12'd3048] = 8'd209;
vramDataLower[12'd3049] = 8'd147;
vramDataLower[12'd3050] = 8'd202;
vramDataLower[12'd3051] = 8'd147;
vramDataLower[12'd3052] = 8'd135;
vramDataLower[12'd3053] = 8'd55;
vramDataLower[12'd3054] = 8'd214;
vramDataLower[12'd3055] = 8'd55;
vramDataLower[12'd3056] = 8'd95;
vramDataLower[12'd3057] = 8'd135;
vramDataLower[12'd3058] = 8'd210;
vramDataLower[12'd3059] = 8'd135;
vramDataLower[12'd3060] = 8'd155;
vramDataLower[12'd3061] = 8'd135;
vramDataLower[12'd3062] = 8'd16;
vramDataLower[12'd3063] = 8'd120;
vramDataLower[12'd3064] = 8'd108;
vramDataLower[12'd3065] = 8'd8;
vramDataLower[12'd3066] = 8'd96;
vramDataLower[12'd3067] = 8'd8;
vramDataLower[12'd3068] = 8'd214;
vramDataLower[12'd3069] = 8'd8;
vramDataLower[12'd3070] = 8'd94;
vramDataLower[12'd3071] = 8'd120;
vramDataLower[12'd3072] = 8'd252;
vramDataLower[12'd3073] = 8'd152;
vramDataLower[12'd3074] = 8'd252;
vramDataLower[12'd3075] = 8'd152;
vramDataLower[12'd3076] = 8'd200;
vramDataLower[12'd3077] = 8'd120;
vramDataLower[12'd3078] = 8'd16;
vramDataLower[12'd3079] = 8'd135;
vramDataLower[12'd3080] = 8'd110;
vramDataLower[12'd3081] = 8'd247;
vramDataLower[12'd3082] = 8'd219;
vramDataLower[12'd3083] = 8'd123;
vramDataLower[12'd3084] = 8'd96;
vramDataLower[12'd3085] = 8'd247;
vramDataLower[12'd3086] = 8'd196;
vramDataLower[12'd3087] = 8'd247;
vramDataLower[12'd3088] = 8'd30;
vramDataLower[12'd3089] = 8'd87;
vramDataLower[12'd3090] = 8'd93;
vramDataLower[12'd3091] = 8'd135;
vramDataLower[12'd3092] = 8'd116;
vramDataLower[12'd3093] = 8'd119;
vramDataLower[12'd3094] = 8'd17;
vramDataLower[12'd3095] = 8'd247;
vramDataLower[12'd3096] = 8'd251;
vramDataLower[12'd3097] = 8'd247;
vramDataLower[12'd3098] = 8'd16;
vramDataLower[12'd3099] = 8'd247;
vramDataLower[12'd3100] = 8'd251;
vramDataLower[12'd3101] = 8'd135;
vramDataLower[12'd3102] = 8'd210;
vramDataLower[12'd3103] = 8'd135;
vramDataLower[12'd3104] = 8'd37;
vramDataLower[12'd3105] = 8'd135;
vramDataLower[12'd3106] = 8'd244;
vramDataLower[12'd3107] = 8'd135;
vramDataLower[12'd3108] = 8'd101;
vramDataLower[12'd3109] = 8'd135;
vramDataLower[12'd3110] = 8'd30;
vramDataLower[12'd3111] = 8'd135;
vramDataLower[12'd3112] = 8'd97;
vramDataLower[12'd3113] = 8'd135;
vramDataLower[12'd3114] = 8'd148;
vramDataLower[12'd3115] = 8'd120;
vramDataLower[12'd3116] = 8'd30;
vramDataLower[12'd3117] = 8'd120;
vramDataLower[12'd3118] = 8'd83;
vramDataLower[12'd3119] = 8'd120;
vramDataLower[12'd3120] = 8'd135;
vramDataLower[12'd3121] = 8'd120;
vramDataLower[12'd3122] = 8'd164;
vramDataLower[12'd3123] = 8'd120;
vramDataLower[12'd3124] = 8'd210;
vramDataLower[12'd3125] = 8'd120;
vramDataLower[12'd3126] = 8'd155;
vramDataLower[12'd3127] = 8'd120;
vramDataLower[12'd3128] = 8'd202;
vramDataLower[12'd3129] = 8'd135;
vramDataLower[12'd3130] = 8'd30;
vramDataLower[12'd3131] = 8'd120;
vramDataLower[12'd3132] = 8'd70;
vramDataLower[12'd3133] = 8'd120;
vramDataLower[12'd3134] = 8'd135;
vramDataLower[12'd3135] = 8'd120;
vramDataLower[12'd3136] = 8'd135;
vramDataLower[12'd3137] = 8'd120;
vramDataLower[12'd3138] = 8'd30;
vramDataLower[12'd3139] = 8'd120;
vramDataLower[12'd3140] = 8'd18;
vramDataLower[12'd3141] = 8'd152;
vramDataLower[12'd3142] = 8'd214;
vramDataLower[12'd3143] = 8'd120;
vramDataLower[12'd3144] = 8'd240;
vramDataLower[12'd3145] = 8'd120;
vramDataLower[12'd3146] = 8'd210;
vramDataLower[12'd3147] = 8'd120;
vramDataLower[12'd3148] = 8'd17;
vramDataLower[12'd3149] = 8'd120;
vramDataLower[12'd3150] = 8'd101;
vramDataLower[12'd3151] = 8'd120;
vramDataLower[12'd3152] = 8'd214;
vramDataLower[12'd3153] = 8'd120;
vramDataLower[12'd3154] = 8'd80;
vramDataLower[12'd3155] = 8'd135;
vramDataLower[12'd3156] = 8'd115;
vramDataLower[12'd3157] = 8'd135;
vramDataLower[12'd3158] = 8'd70;
vramDataLower[12'd3159] = 8'd135;
vramDataLower[12'd3160] = 8'd31;
vramDataLower[12'd3161] = 8'd135;
vramDataLower[12'd3162] = 8'd31;
vramDataLower[12'd3163] = 8'd135;
vramDataLower[12'd3164] = 8'd94;
vramDataLower[12'd3165] = 8'd135;
vramDataLower[12'd3166] = 8'd248;
vramDataLower[12'd3167] = 8'd135;
vramDataLower[12'd3168] = 8'd92;
vramDataLower[12'd3169] = 8'd135;
vramDataLower[12'd3170] = 8'd83;
vramDataLower[12'd3171] = 8'd135;
vramDataLower[12'd3172] = 8'd200;
vramDataLower[12'd3173] = 8'd135;
vramDataLower[12'd3174] = 8'd80;
vramDataLower[12'd3175] = 8'd87;
vramDataLower[12'd3176] = 8'd184;
vramDataLower[12'd3177] = 8'd135;
vramDataLower[12'd3178] = 8'd28;
vramDataLower[12'd3179] = 8'd87;
vramDataLower[12'd3180] = 8'd29;
vramDataLower[12'd3181] = 8'd247;
vramDataLower[12'd3182] = 8'd95;
vramDataLower[12'd3183] = 8'd247;
vramDataLower[12'd3184] = 8'd200;
vramDataLower[12'd3185] = 8'd247;
vramDataLower[12'd3186] = 8'd16;
vramDataLower[12'd3187] = 8'd247;
vramDataLower[12'd3188] = 8'd198;
vramDataLower[12'd3189] = 8'd55;
vramDataLower[12'd3190] = 8'd16;
vramDataLower[12'd3191] = 8'd115;
vramDataLower[12'd3192] = 8'd210;
vramDataLower[12'd3193] = 8'd115;
vramDataLower[12'd3194] = 8'd202;
vramDataLower[12'd3195] = 8'd147;
vramDataLower[12'd3196] = 8'd202;
vramDataLower[12'd3197] = 8'd19;
vramDataLower[12'd3198] = 8'd210;
vramDataLower[12'd3199] = 8'd49;
vramDataLower[12'd3200] = 8'd202;
vramDataLower[12'd3201] = 8'd56;
vramDataLower[12'd3202] = 8'd210;
vramDataLower[12'd3203] = 8'd131;
vramDataLower[12'd3204] = 8'd202;
vramDataLower[12'd3205] = 8'd147;
vramDataLower[12'd3206] = 8'd202;
vramDataLower[12'd3207] = 8'd147;
vramDataLower[12'd3208] = 8'd202;
vramDataLower[12'd3209] = 8'd147;
vramDataLower[12'd3210] = 8'd80;
vramDataLower[12'd3211] = 8'd147;
vramDataLower[12'd3212] = 8'd80;
vramDataLower[12'd3213] = 8'd147;
vramDataLower[12'd3214] = 8'd16;
vramDataLower[12'd3215] = 8'd55;
vramDataLower[12'd3216] = 8'd80;
vramDataLower[12'd3217] = 8'd135;
vramDataLower[12'd3218] = 8'd226;
vramDataLower[12'd3219] = 8'd135;
vramDataLower[12'd3220] = 8'd228;
vramDataLower[12'd3221] = 8'd135;
vramDataLower[12'd3222] = 8'd0;
vramDataLower[12'd3223] = 8'd199;
vramDataLower[12'd3224] = 8'd16;
vramDataLower[12'd3225] = 8'd120;
vramDataLower[12'd3226] = 8'd209;
vramDataLower[12'd3227] = 8'd8;
vramDataLower[12'd3228] = 8'd16;
vramDataLower[12'd3229] = 8'd8;
vramDataLower[12'd3230] = 8'd81;
vramDataLower[12'd3231] = 8'd136;
vramDataLower[12'd3232] = 8'd95;
vramDataLower[12'd3233] = 8'd8;
vramDataLower[12'd3234] = 8'd183;
vramDataLower[12'd3235] = 8'd8;
vramDataLower[12'd3236] = 8'd95;
vramDataLower[12'd3237] = 8'd8;
vramDataLower[12'd3238] = 8'd94;
vramDataLower[12'd3239] = 8'd120;
vramDataLower[12'd3240] = 8'd223;
vramDataLower[12'd3241] = 8'd120;
vramDataLower[12'd3242] = 8'd223;
vramDataLower[12'd3243] = 8'd120;
vramDataLower[12'd3244] = 8'd183;
vramDataLower[12'd3245] = 8'd135;
vramDataLower[12'd3246] = 8'd210;
vramDataLower[12'd3247] = 8'd135;
vramDataLower[12'd3248] = 8'd230;
vramDataLower[12'd3249] = 8'd135;
vramDataLower[12'd3250] = 8'd31;
vramDataLower[12'd3251] = 8'd247;
vramDataLower[12'd3252] = 8'd208;
vramDataLower[12'd3253] = 8'd247;
vramDataLower[12'd3254] = 8'd248;
vramDataLower[12'd3255] = 8'd247;
vramDataLower[12'd3256] = 8'd200;
vramDataLower[12'd3257] = 8'd247;
vramDataLower[12'd3258] = 8'd155;
vramDataLower[12'd3259] = 8'd247;
vramDataLower[12'd3260] = 8'd28;
vramDataLower[12'd3261] = 8'd247;
vramDataLower[12'd3262] = 8'd155;
vramDataLower[12'd3263] = 8'd135;
vramDataLower[12'd3264] = 8'd149;
vramDataLower[12'd3265] = 8'd135;
vramDataLower[12'd3266] = 8'd240;
vramDataLower[12'd3267] = 8'd135;
vramDataLower[12'd3268] = 8'd31;
vramDataLower[12'd3269] = 8'd135;
vramDataLower[12'd3270] = 8'd101;
vramDataLower[12'd3271] = 8'd120;
vramDataLower[12'd3272] = 8'd135;
vramDataLower[12'd3273] = 8'd135;
vramDataLower[12'd3274] = 8'd90;
vramDataLower[12'd3275] = 8'd135;
vramDataLower[12'd3276] = 8'd156;
vramDataLower[12'd3277] = 8'd135;
vramDataLower[12'd3278] = 8'd155;
vramDataLower[12'd3279] = 8'd120;
vramDataLower[12'd3280] = 8'd37;
vramDataLower[12'd3281] = 8'd120;
vramDataLower[12'd3282] = 8'd156;
vramDataLower[12'd3283] = 8'd120;
vramDataLower[12'd3284] = 8'd202;
vramDataLower[12'd3285] = 8'd120;
vramDataLower[12'd3286] = 8'd83;
vramDataLower[12'd3287] = 8'd120;
vramDataLower[12'd3288] = 8'd17;
vramDataLower[12'd3289] = 8'd120;
vramDataLower[12'd3290] = 8'd145;
vramDataLower[12'd3291] = 8'd120;
vramDataLower[12'd3292] = 8'd30;
vramDataLower[12'd3293] = 8'd120;
vramDataLower[12'd3294] = 8'd101;
vramDataLower[12'd3295] = 8'd120;
vramDataLower[12'd3296] = 8'd202;
vramDataLower[12'd3297] = 8'd120;
vramDataLower[12'd3298] = 8'd30;
vramDataLower[12'd3299] = 8'd120;
vramDataLower[12'd3300] = 8'd83;
vramDataLower[12'd3301] = 8'd120;
vramDataLower[12'd3302] = 8'd83;
vramDataLower[12'd3303] = 8'd120;
vramDataLower[12'd3304] = 8'd30;
vramDataLower[12'd3305] = 8'd120;
vramDataLower[12'd3306] = 8'd80;
vramDataLower[12'd3307] = 8'd135;
vramDataLower[12'd3308] = 8'd80;
vramDataLower[12'd3309] = 8'd120;
vramDataLower[12'd3310] = 8'd164;
vramDataLower[12'd3311] = 8'd135;
vramDataLower[12'd3312] = 8'd31;
vramDataLower[12'd3313] = 8'd135;
vramDataLower[12'd3314] = 8'd16;
vramDataLower[12'd3315] = 8'd135;
vramDataLower[12'd3316] = 8'd200;
vramDataLower[12'd3317] = 8'd135;
vramDataLower[12'd3318] = 8'd17;
vramDataLower[12'd3319] = 8'd135;
vramDataLower[12'd3320] = 8'd248;
vramDataLower[12'd3321] = 8'd135;
vramDataLower[12'd3322] = 8'd253;
vramDataLower[12'd3323] = 8'd103;
vramDataLower[12'd3324] = 8'd150;
vramDataLower[12'd3325] = 8'd119;
vramDataLower[12'd3326] = 8'd251;
vramDataLower[12'd3327] = 8'd55;
vramDataLower[12'd3328] = 8'd83;
vramDataLower[12'd3329] = 8'd135;
vramDataLower[12'd3330] = 8'd249;
vramDataLower[12'd3331] = 8'd135;
vramDataLower[12'd3332] = 8'd31;
vramDataLower[12'd3333] = 8'd135;
vramDataLower[12'd3334] = 8'd31;
vramDataLower[12'd3335] = 8'd135;
vramDataLower[12'd3336] = 8'd191;
vramDataLower[12'd3337] = 8'd135;
vramDataLower[12'd3338] = 8'd170;
vramDataLower[12'd3339] = 8'd247;
vramDataLower[12'd3340] = 8'd95;
vramDataLower[12'd3341] = 8'd247;
vramDataLower[12'd3342] = 8'd198;
vramDataLower[12'd3343] = 8'd247;
vramDataLower[12'd3344] = 8'd202;
vramDataLower[12'd3345] = 8'd247;
vramDataLower[12'd3346] = 8'd16;
vramDataLower[12'd3347] = 8'd247;
vramDataLower[12'd3348] = 8'd80;
vramDataLower[12'd3349] = 8'd115;
vramDataLower[12'd3350] = 8'd31;
vramDataLower[12'd3351] = 8'd147;
vramDataLower[12'd3352] = 8'd16;
vramDataLower[12'd3353] = 8'd147;
vramDataLower[12'd3354] = 8'd210;
vramDataLower[12'd3355] = 8'd19;
vramDataLower[12'd3356] = 8'd210;
vramDataLower[12'd3357] = 8'd131;
vramDataLower[12'd3358] = 8'd210;
vramDataLower[12'd3359] = 8'd131;
vramDataLower[12'd3360] = 8'd202;
vramDataLower[12'd3361] = 8'd24;
vramDataLower[12'd3362] = 8'd202;
vramDataLower[12'd3363] = 8'd56;
vramDataLower[12'd3364] = 8'd145;
vramDataLower[12'd3365] = 8'd56;
vramDataLower[12'd3366] = 8'd16;
vramDataLower[12'd3367] = 8'd56;
vramDataLower[12'd3368] = 8'd202;
vramDataLower[12'd3369] = 8'd24;
vramDataLower[12'd3370] = 8'd37;
vramDataLower[12'd3371] = 8'd8;
vramDataLower[12'd3372] = 8'd16;
vramDataLower[12'd3373] = 8'd8;
vramDataLower[12'd3374] = 8'd198;
vramDataLower[12'd3375] = 8'd152;
vramDataLower[12'd3376] = 8'd37;
vramDataLower[12'd3377] = 8'd135;
vramDataLower[12'd3378] = 8'd16;
vramDataLower[12'd3379] = 8'd135;
vramDataLower[12'd3380] = 8'd16;
vramDataLower[12'd3381] = 8'd135;
vramDataLower[12'd3382] = 8'd166;
vramDataLower[12'd3383] = 8'd87;
vramDataLower[12'd3384] = 8'd221;
vramDataLower[12'd3385] = 8'd120;
vramDataLower[12'd3386] = 8'd202;
vramDataLower[12'd3387] = 8'd8;
vramDataLower[12'd3388] = 8'd16;
vramDataLower[12'd3389] = 8'd8;
vramDataLower[12'd3390] = 8'd52;
vramDataLower[12'd3391] = 8'd200;
vramDataLower[12'd3392] = 8'd168;
vramDataLower[12'd3393] = 8'd120;
vramDataLower[12'd3394] = 8'd198;
vramDataLower[12'd3395] = 8'd8;
vramDataLower[12'd3396] = 8'd80;
vramDataLower[12'd3397] = 8'd8;
vramDataLower[12'd3398] = 8'd95;
vramDataLower[12'd3399] = 8'd120;
vramDataLower[12'd3400] = 8'd214;
vramDataLower[12'd3401] = 8'd120;
vramDataLower[12'd3402] = 8'd214;
vramDataLower[12'd3403] = 8'd120;
vramDataLower[12'd3404] = 8'd223;
vramDataLower[12'd3405] = 8'd135;
vramDataLower[12'd3406] = 8'd252;
vramDataLower[12'd3407] = 8'd135;
vramDataLower[12'd3408] = 8'd60;
vramDataLower[12'd3409] = 8'd247;
vramDataLower[12'd3410] = 8'd243;
vramDataLower[12'd3411] = 8'd247;
vramDataLower[12'd3412] = 8'd18;
vramDataLower[12'd3413] = 8'd247;
vramDataLower[12'd3414] = 8'd240;
vramDataLower[12'd3415] = 8'd247;
vramDataLower[12'd3416] = 8'd212;
vramDataLower[12'd3417] = 8'd247;
vramDataLower[12'd3418] = 8'd166;
vramDataLower[12'd3419] = 8'd135;
vramDataLower[12'd3420] = 8'd210;
vramDataLower[12'd3421] = 8'd135;
vramDataLower[12'd3422] = 8'd135;
vramDataLower[12'd3423] = 8'd135;
vramDataLower[12'd3424] = 8'd67;
vramDataLower[12'd3425] = 8'd135;
vramDataLower[12'd3426] = 8'd122;
vramDataLower[12'd3427] = 8'd135;
vramDataLower[12'd3428] = 8'd209;
vramDataLower[12'd3429] = 8'd135;
vramDataLower[12'd3430] = 8'd83;
vramDataLower[12'd3431] = 8'd135;
vramDataLower[12'd3432] = 8'd228;
vramDataLower[12'd3433] = 8'd120;
vramDataLower[12'd3434] = 8'd31;
vramDataLower[12'd3435] = 8'd135;
vramDataLower[12'd3436] = 8'd202;
vramDataLower[12'd3437] = 8'd135;
vramDataLower[12'd3438] = 8'd31;
vramDataLower[12'd3439] = 8'd135;
vramDataLower[12'd3440] = 8'd80;
vramDataLower[12'd3441] = 8'd120;
vramDataLower[12'd3442] = 8'd208;
vramDataLower[12'd3443] = 8'd120;
vramDataLower[12'd3444] = 8'd240;
vramDataLower[12'd3445] = 8'd120;
vramDataLower[12'd3446] = 8'd205;
vramDataLower[12'd3447] = 8'd120;
vramDataLower[12'd3448] = 8'd239;
vramDataLower[12'd3449] = 8'd120;
vramDataLower[12'd3450] = 8'd31;
vramDataLower[12'd3451] = 8'd120;
vramDataLower[12'd3452] = 8'd30;
vramDataLower[12'd3453] = 8'd120;
vramDataLower[12'd3454] = 8'd31;
vramDataLower[12'd3455] = 8'd120;
vramDataLower[12'd3456] = 8'd31;
vramDataLower[12'd3457] = 8'd120;
vramDataLower[12'd3458] = 8'd239;
vramDataLower[12'd3459] = 8'd120;
vramDataLower[12'd3460] = 8'd83;
vramDataLower[12'd3461] = 8'd120;
vramDataLower[12'd3462] = 8'd37;
vramDataLower[12'd3463] = 8'd120;
vramDataLower[12'd3464] = 8'd240;
vramDataLower[12'd3465] = 8'd135;
vramDataLower[12'd3466] = 8'd31;
vramDataLower[12'd3467] = 8'd135;
vramDataLower[12'd3468] = 8'd30;
vramDataLower[12'd3469] = 8'd135;
vramDataLower[12'd3470] = 8'd145;
vramDataLower[12'd3471] = 8'd135;
vramDataLower[12'd3472] = 8'd156;
vramDataLower[12'd3473] = 8'd135;
vramDataLower[12'd3474] = 8'd90;
vramDataLower[12'd3475] = 8'd135;
vramDataLower[12'd3476] = 8'd95;
vramDataLower[12'd3477] = 8'd135;
vramDataLower[12'd3478] = 8'd115;
vramDataLower[12'd3479] = 8'd135;
vramDataLower[12'd3480] = 8'd67;
vramDataLower[12'd3481] = 8'd135;
vramDataLower[12'd3482] = 8'd228;
vramDataLower[12'd3483] = 8'd135;
vramDataLower[12'd3484] = 8'd95;
vramDataLower[12'd3485] = 8'd135;
vramDataLower[12'd3486] = 8'd31;
vramDataLower[12'd3487] = 8'd135;
vramDataLower[12'd3488] = 8'd29;
vramDataLower[12'd3489] = 8'd135;
vramDataLower[12'd3490] = 8'd135;
vramDataLower[12'd3491] = 8'd135;
vramDataLower[12'd3492] = 8'd190;
vramDataLower[12'd3493] = 8'd135;
vramDataLower[12'd3494] = 8'd211;
vramDataLower[12'd3495] = 8'd135;
vramDataLower[12'd3496] = 8'd248;
vramDataLower[12'd3497] = 8'd135;
vramDataLower[12'd3498] = 8'd170;
vramDataLower[12'd3499] = 8'd247;
vramDataLower[12'd3500] = 8'd50;
vramDataLower[12'd3501] = 8'd247;
vramDataLower[12'd3502] = 8'd30;
vramDataLower[12'd3503] = 8'd247;
vramDataLower[12'd3504] = 8'd210;
vramDataLower[12'd3505] = 8'd247;
vramDataLower[12'd3506] = 8'd16;
vramDataLower[12'd3507] = 8'd247;
vramDataLower[12'd3508] = 8'd16;
vramDataLower[12'd3509] = 8'd115;
vramDataLower[12'd3510] = 8'd210;
vramDataLower[12'd3511] = 8'd131;
vramDataLower[12'd3512] = 8'd210;
vramDataLower[12'd3513] = 8'd131;
vramDataLower[12'd3514] = 8'd202;
vramDataLower[12'd3515] = 8'd56;
vramDataLower[12'd3516] = 8'd209;
vramDataLower[12'd3517] = 8'd56;
vramDataLower[12'd3518] = 8'd209;
vramDataLower[12'd3519] = 8'd56;
vramDataLower[12'd3520] = 8'd210;
vramDataLower[12'd3521] = 8'd24;
vramDataLower[12'd3522] = 8'd210;
vramDataLower[12'd3523] = 8'd24;
vramDataLower[12'd3524] = 8'd202;
vramDataLower[12'd3525] = 8'd56;
vramDataLower[12'd3526] = 8'd148;
vramDataLower[12'd3527] = 8'd56;
vramDataLower[12'd3528] = 8'd16;
vramDataLower[12'd3529] = 8'd56;
vramDataLower[12'd3530] = 8'd127;
vramDataLower[12'd3531] = 8'd120;
vramDataLower[12'd3532] = 8'd30;
vramDataLower[12'd3533] = 8'd120;
vramDataLower[12'd3534] = 8'd31;
vramDataLower[12'd3535] = 8'd120;
vramDataLower[12'd3536] = 8'd200;
vramDataLower[12'd3537] = 8'd120;
vramDataLower[12'd3538] = 8'd210;
vramDataLower[12'd3539] = 8'd135;
vramDataLower[12'd3540] = 8'd210;
vramDataLower[12'd3541] = 8'd135;
vramDataLower[12'd3542] = 8'd16;
vramDataLower[12'd3543] = 8'd135;
vramDataLower[12'd3544] = 8'd212;
vramDataLower[12'd3545] = 8'd55;
vramDataLower[12'd3546] = 8'd16;
vramDataLower[12'd3547] = 8'd120;
vramDataLower[12'd3548] = 8'd83;
vramDataLower[12'd3549] = 8'd8;
vramDataLower[12'd3550] = 8'd80;
vramDataLower[12'd3551] = 8'd8;
vramDataLower[12'd3552] = 8'd16;
vramDataLower[12'd3553] = 8'd8;
vramDataLower[12'd3554] = 8'd172;
vramDataLower[12'd3555] = 8'd120;
vramDataLower[12'd3556] = 8'd164;
vramDataLower[12'd3557] = 8'd135;
vramDataLower[12'd3558] = 8'd94;
vramDataLower[12'd3559] = 8'd135;
vramDataLower[12'd3560] = 8'd141;
vramDataLower[12'd3561] = 8'd135;
vramDataLower[12'd3562] = 8'd145;
vramDataLower[12'd3563] = 8'd247;
vramDataLower[12'd3564] = 8'd139;
vramDataLower[12'd3565] = 8'd247;
vramDataLower[12'd3566] = 8'd211;
vramDataLower[12'd3567] = 8'd247;
vramDataLower[12'd3568] = 8'd45;
vramDataLower[12'd3569] = 8'd135;
vramDataLower[12'd3570] = 8'd46;
vramDataLower[12'd3571] = 8'd135;
vramDataLower[12'd3572] = 8'd192;
vramDataLower[12'd3573] = 8'd247;
vramDataLower[12'd3574] = 8'd92;
vramDataLower[12'd3575] = 8'd135;
vramDataLower[12'd3576] = 8'd127;
vramDataLower[12'd3577] = 8'd135;
vramDataLower[12'd3578] = 8'd218;
vramDataLower[12'd3579] = 8'd135;
vramDataLower[12'd3580] = 8'd200;
vramDataLower[12'd3581] = 8'd135;
vramDataLower[12'd3582] = 8'd240;
vramDataLower[12'd3583] = 8'd135;
vramDataLower[12'd3584] = 8'd9;
vramDataLower[12'd3585] = 8'd135;
vramDataLower[12'd3586] = 8'd230;
vramDataLower[12'd3587] = 8'd135;
vramDataLower[12'd3588] = 8'd164;
vramDataLower[12'd3589] = 8'd135;
vramDataLower[12'd3590] = 8'd240;
vramDataLower[12'd3591] = 8'd120;
vramDataLower[12'd3592] = 8'd83;
vramDataLower[12'd3593] = 8'd120;
vramDataLower[12'd3594] = 8'd90;
vramDataLower[12'd3595] = 8'd120;
vramDataLower[12'd3596] = 8'd42;
vramDataLower[12'd3597] = 8'd120;
vramDataLower[12'd3598] = 8'd16;
vramDataLower[12'd3599] = 8'd135;
vramDataLower[12'd3600] = 8'd240;
vramDataLower[12'd3601] = 8'd120;
vramDataLower[12'd3602] = 8'd30;
vramDataLower[12'd3603] = 8'd135;
vramDataLower[12'd3604] = 8'd115;
vramDataLower[12'd3605] = 8'd120;
vramDataLower[12'd3606] = 8'd122;
vramDataLower[12'd3607] = 8'd120;
vramDataLower[12'd3608] = 8'd240;
vramDataLower[12'd3609] = 8'd120;
vramDataLower[12'd3610] = 8'd31;
vramDataLower[12'd3611] = 8'd120;
vramDataLower[12'd3612] = 8'd30;
vramDataLower[12'd3613] = 8'd120;
vramDataLower[12'd3614] = 8'd83;
vramDataLower[12'd3615] = 8'd120;
vramDataLower[12'd3616] = 8'd155;
vramDataLower[12'd3617] = 8'd120;
vramDataLower[12'd3618] = 8'd211;
vramDataLower[12'd3619] = 8'd120;
vramDataLower[12'd3620] = 8'd83;
vramDataLower[12'd3621] = 8'd120;
vramDataLower[12'd3622] = 8'd80;
vramDataLower[12'd3623] = 8'd135;
vramDataLower[12'd3624] = 8'd80;
vramDataLower[12'd3625] = 8'd135;
vramDataLower[12'd3626] = 8'd30;
vramDataLower[12'd3627] = 8'd135;
vramDataLower[12'd3628] = 8'd90;
vramDataLower[12'd3629] = 8'd135;
vramDataLower[12'd3630] = 8'd210;
vramDataLower[12'd3631] = 8'd135;
vramDataLower[12'd3632] = 8'd50;
vramDataLower[12'd3633] = 8'd135;
vramDataLower[12'd3634] = 8'd37;
vramDataLower[12'd3635] = 8'd135;
vramDataLower[12'd3636] = 8'd135;
vramDataLower[12'd3637] = 8'd135;
vramDataLower[12'd3638] = 8'd31;
vramDataLower[12'd3639] = 8'd135;
vramDataLower[12'd3640] = 8'd251;
vramDataLower[12'd3641] = 8'd135;
vramDataLower[12'd3642] = 8'd90;
vramDataLower[12'd3643] = 8'd135;
vramDataLower[12'd3644] = 8'd30;
vramDataLower[12'd3645] = 8'd135;
vramDataLower[12'd3646] = 8'd228;
vramDataLower[12'd3647] = 8'd55;
vramDataLower[12'd3648] = 8'd248;
vramDataLower[12'd3649] = 8'd135;
vramDataLower[12'd3650] = 8'd207;
vramDataLower[12'd3651] = 8'd135;
vramDataLower[12'd3652] = 8'd51;
vramDataLower[12'd3653] = 8'd135;
vramDataLower[12'd3654] = 8'd28;
vramDataLower[12'd3655] = 8'd135;
vramDataLower[12'd3656] = 8'd96;
vramDataLower[12'd3657] = 8'd135;
vramDataLower[12'd3658] = 8'd95;
vramDataLower[12'd3659] = 8'd247;
vramDataLower[12'd3660] = 8'd30;
vramDataLower[12'd3661] = 8'd247;
vramDataLower[12'd3662] = 8'd148;
vramDataLower[12'd3663] = 8'd247;
vramDataLower[12'd3664] = 8'd16;
vramDataLower[12'd3665] = 8'd247;
vramDataLower[12'd3666] = 8'd198;
vramDataLower[12'd3667] = 8'd55;
vramDataLower[12'd3668] = 8'd16;
vramDataLower[12'd3669] = 8'd115;
vramDataLower[12'd3670] = 8'd210;
vramDataLower[12'd3671] = 8'd147;
vramDataLower[12'd3672] = 8'd210;
vramDataLower[12'd3673] = 8'd147;
vramDataLower[12'd3674] = 8'd202;
vramDataLower[12'd3675] = 8'd19;
vramDataLower[12'd3676] = 8'd202;
vramDataLower[12'd3677] = 8'd19;
vramDataLower[12'd3678] = 8'd202;
vramDataLower[12'd3679] = 8'd19;
vramDataLower[12'd3680] = 8'd202;
vramDataLower[12'd3681] = 8'd24;
vramDataLower[12'd3682] = 8'd202;
vramDataLower[12'd3683] = 8'd24;
vramDataLower[12'd3684] = 8'd202;
vramDataLower[12'd3685] = 8'd152;
vramDataLower[12'd3686] = 8'd202;
vramDataLower[12'd3687] = 8'd56;
vramDataLower[12'd3688] = 8'd202;
vramDataLower[12'd3689] = 8'd152;
vramDataLower[12'd3690] = 8'd210;
vramDataLower[12'd3691] = 8'd152;
vramDataLower[12'd3692] = 8'd210;
vramDataLower[12'd3693] = 8'd152;
vramDataLower[12'd3694] = 8'd135;
vramDataLower[12'd3695] = 8'd152;
vramDataLower[12'd3696] = 8'd214;
vramDataLower[12'd3697] = 8'd152;
vramDataLower[12'd3698] = 8'd210;
vramDataLower[12'd3699] = 8'd120;
vramDataLower[12'd3700] = 8'd209;
vramDataLower[12'd3701] = 8'd120;
vramDataLower[12'd3702] = 8'd80;
vramDataLower[12'd3703] = 8'd135;
vramDataLower[12'd3704] = 8'd214;
vramDataLower[12'd3705] = 8'd135;
vramDataLower[12'd3706] = 8'd16;
vramDataLower[12'd3707] = 8'd120;
vramDataLower[12'd3708] = 8'd117;
vramDataLower[12'd3709] = 8'd152;
vramDataLower[12'd3710] = 8'd45;
vramDataLower[12'd3711] = 8'd8;
vramDataLower[12'd3712] = 8'd88;
vramDataLower[12'd3713] = 8'd120;
vramDataLower[12'd3714] = 8'd95;
vramDataLower[12'd3715] = 8'd135;
vramDataLower[12'd3716] = 8'd252;
vramDataLower[12'd3717] = 8'd135;
vramDataLower[12'd3718] = 8'd247;
vramDataLower[12'd3719] = 8'd247;
vramDataLower[12'd3720] = 8'd94;
vramDataLower[12'd3721] = 8'd135;
vramDataLower[12'd3722] = 8'd62;
vramDataLower[12'd3723] = 8'd135;
vramDataLower[12'd3724] = 8'd46;
vramDataLower[12'd3725] = 8'd135;
vramDataLower[12'd3726] = 8'd252;
vramDataLower[12'd3727] = 8'd135;
vramDataLower[12'd3728] = 8'd96;
vramDataLower[12'd3729] = 8'd247;
vramDataLower[12'd3730] = 8'd30;
vramDataLower[12'd3731] = 8'd135;
vramDataLower[12'd3732] = 8'd16;
vramDataLower[12'd3733] = 8'd135;
vramDataLower[12'd3734] = 8'd149;
vramDataLower[12'd3735] = 8'd135;
vramDataLower[12'd3736] = 8'd171;
vramDataLower[12'd3737] = 8'd120;
vramDataLower[12'd3738] = 8'd51;
vramDataLower[12'd3739] = 8'd120;
vramDataLower[12'd3740] = 8'd85;
vramDataLower[12'd3741] = 8'd135;
vramDataLower[12'd3742] = 8'd200;
vramDataLower[12'd3743] = 8'd120;
vramDataLower[12'd3744] = 8'd83;
vramDataLower[12'd3745] = 8'd135;
vramDataLower[12'd3746] = 8'd55;
vramDataLower[12'd3747] = 8'd135;
vramDataLower[12'd3748] = 8'd9;
vramDataLower[12'd3749] = 8'd120;
vramDataLower[12'd3750] = 8'd164;
vramDataLower[12'd3751] = 8'd135;
vramDataLower[12'd3752] = 8'd83;
vramDataLower[12'd3753] = 8'd120;
vramDataLower[12'd3754] = 8'd166;
vramDataLower[12'd3755] = 8'd120;
vramDataLower[12'd3756] = 8'd31;
vramDataLower[12'd3757] = 8'd120;
vramDataLower[12'd3758] = 8'd115;
vramDataLower[12'd3759] = 8'd120;
vramDataLower[12'd3760] = 8'd16;
vramDataLower[12'd3761] = 8'd135;
vramDataLower[12'd3762] = 8'd171;
vramDataLower[12'd3763] = 8'd135;
vramDataLower[12'd3764] = 8'd208;
vramDataLower[12'd3765] = 8'd135;
vramDataLower[12'd3766] = 8'd31;
vramDataLower[12'd3767] = 8'd120;
vramDataLower[12'd3768] = 8'd145;
vramDataLower[12'd3769] = 8'd120;
vramDataLower[12'd3770] = 8'd30;
vramDataLower[12'd3771] = 8'd120;
vramDataLower[12'd3772] = 8'd135;
vramDataLower[12'd3773] = 8'd120;
vramDataLower[12'd3774] = 8'd16;
vramDataLower[12'd3775] = 8'd120;
vramDataLower[12'd3776] = 8'd135;
vramDataLower[12'd3777] = 8'd120;
vramDataLower[12'd3778] = 8'd210;
vramDataLower[12'd3779] = 8'd120;
vramDataLower[12'd3780] = 8'd31;
vramDataLower[12'd3781] = 8'd135;
vramDataLower[12'd3782] = 8'd148;
vramDataLower[12'd3783] = 8'd120;
vramDataLower[12'd3784] = 8'd164;
vramDataLower[12'd3785] = 8'd120;
vramDataLower[12'd3786] = 8'd80;
vramDataLower[12'd3787] = 8'd120;
vramDataLower[12'd3788] = 8'd228;
vramDataLower[12'd3789] = 8'd120;
vramDataLower[12'd3790] = 8'd200;
vramDataLower[12'd3791] = 8'd120;
vramDataLower[12'd3792] = 8'd145;
vramDataLower[12'd3793] = 8'd135;
vramDataLower[12'd3794] = 8'd95;
vramDataLower[12'd3795] = 8'd135;
vramDataLower[12'd3796] = 8'd90;
vramDataLower[12'd3797] = 8'd135;
vramDataLower[12'd3798] = 8'd210;
vramDataLower[12'd3799] = 8'd135;
vramDataLower[12'd3800] = 8'd238;
vramDataLower[12'd3801] = 8'd135;
vramDataLower[12'd3802] = 8'd91;
vramDataLower[12'd3803] = 8'd135;
vramDataLower[12'd3804] = 8'd240;
vramDataLower[12'd3805] = 8'd135;
vramDataLower[12'd3806] = 8'd229;
vramDataLower[12'd3807] = 8'd55;
vramDataLower[12'd3808] = 8'd90;
vramDataLower[12'd3809] = 8'd55;
vramDataLower[12'd3810] = 8'd250;
vramDataLower[12'd3811] = 8'd135;
vramDataLower[12'd3812] = 8'd30;
vramDataLower[12'd3813] = 8'd135;
vramDataLower[12'd3814] = 8'd228;
vramDataLower[12'd3815] = 8'd135;
vramDataLower[12'd3816] = 8'd116;
vramDataLower[12'd3817] = 8'd87;
vramDataLower[12'd3818] = 8'd148;
vramDataLower[12'd3819] = 8'd119;
vramDataLower[12'd3820] = 8'd95;
vramDataLower[12'd3821] = 8'd247;
vramDataLower[12'd3822] = 8'd80;
vramDataLower[12'd3823] = 8'd247;
vramDataLower[12'd3824] = 8'd235;
vramDataLower[12'd3825] = 8'd119;
vramDataLower[12'd3826] = 8'd198;
vramDataLower[12'd3827] = 8'd183;
vramDataLower[12'd3828] = 8'd80;
vramDataLower[12'd3829] = 8'd123;
vramDataLower[12'd3830] = 8'd210;
vramDataLower[12'd3831] = 8'd179;
vramDataLower[12'd3832] = 8'd210;
vramDataLower[12'd3833] = 8'd179;
vramDataLower[12'd3834] = 8'd210;
vramDataLower[12'd3835] = 8'd179;
vramDataLower[12'd3836] = 8'd210;
vramDataLower[12'd3837] = 8'd179;
vramDataLower[12'd3838] = 8'd210;
vramDataLower[12'd3839] = 8'd147;
vramDataLower[12'd3840] = 8'd209;
vramDataLower[12'd3841] = 8'd152;
vramDataLower[12'd3842] = 8'd164;
vramDataLower[12'd3843] = 8'd152;
vramDataLower[12'd3844] = 8'd83;
vramDataLower[12'd3845] = 8'd152;
vramDataLower[12'd3846] = 8'd30;
vramDataLower[12'd3847] = 8'd152;
vramDataLower[12'd3848] = 8'd181;
vramDataLower[12'd3849] = 8'd152;
vramDataLower[12'd3850] = 8'd145;
vramDataLower[12'd3851] = 8'd152;
vramDataLower[12'd3852] = 8'd210;
vramDataLower[12'd3853] = 8'd152;
vramDataLower[12'd3854] = 8'd148;
vramDataLower[12'd3855] = 8'd152;
vramDataLower[12'd3856] = 8'd31;
vramDataLower[12'd3857] = 8'd120;
vramDataLower[12'd3858] = 8'd80;
vramDataLower[12'd3859] = 8'd120;
vramDataLower[12'd3860] = 8'd210;
vramDataLower[12'd3861] = 8'd152;
vramDataLower[12'd3862] = 8'd202;
vramDataLower[12'd3863] = 8'd120;
vramDataLower[12'd3864] = 8'd210;
vramDataLower[12'd3865] = 8'd135;
vramDataLower[12'd3866] = 8'd202;
vramDataLower[12'd3867] = 8'd120;
vramDataLower[12'd3868] = 8'd31;
vramDataLower[12'd3869] = 8'd152;
vramDataLower[12'd3870] = 8'd16;
vramDataLower[12'd3871] = 8'd152;
vramDataLower[12'd3872] = 8'd104;
vramDataLower[12'd3873] = 8'd120;
vramDataLower[12'd3874] = 8'd164;
vramDataLower[12'd3875] = 8'd120;
vramDataLower[12'd3876] = 8'd198;
vramDataLower[12'd3877] = 8'd120;
vramDataLower[12'd3878] = 8'd135;
vramDataLower[12'd3879] = 8'd135;
vramDataLower[12'd3880] = 8'd244;
vramDataLower[12'd3881] = 8'd135;
vramDataLower[12'd3882] = 8'd107;
vramDataLower[12'd3883] = 8'd135;
vramDataLower[12'd3884] = 8'd230;
vramDataLower[12'd3885] = 8'd135;
vramDataLower[12'd3886] = 8'd200;
vramDataLower[12'd3887] = 8'd135;
vramDataLower[12'd3888] = 8'd248;
vramDataLower[12'd3889] = 8'd120;
vramDataLower[12'd3890] = 8'd16;
vramDataLower[12'd3891] = 8'd135;
vramDataLower[12'd3892] = 8'd80;
vramDataLower[12'd3893] = 8'd120;
vramDataLower[12'd3894] = 8'd202;
vramDataLower[12'd3895] = 8'd120;
vramDataLower[12'd3896] = 8'd183;
vramDataLower[12'd3897] = 8'd135;
vramDataLower[12'd3898] = 8'd80;
vramDataLower[12'd3899] = 8'd135;
vramDataLower[12'd3900] = 8'd17;
vramDataLower[12'd3901] = 8'd135;
vramDataLower[12'd3902] = 8'd31;
vramDataLower[12'd3903] = 8'd120;
vramDataLower[12'd3904] = 8'd17;
vramDataLower[12'd3905] = 8'd135;
vramDataLower[12'd3906] = 8'd31;
vramDataLower[12'd3907] = 8'd120;
vramDataLower[12'd3908] = 8'd17;
vramDataLower[12'd3909] = 8'd120;
vramDataLower[12'd3910] = 8'd214;
vramDataLower[12'd3911] = 8'd120;
vramDataLower[12'd3912] = 8'd30;
vramDataLower[12'd3913] = 8'd135;
vramDataLower[12'd3914] = 8'd16;
vramDataLower[12'd3915] = 8'd120;
vramDataLower[12'd3916] = 8'd210;
vramDataLower[12'd3917] = 8'd120;
vramDataLower[12'd3918] = 8'd148;
vramDataLower[12'd3919] = 8'd135;
vramDataLower[12'd3920] = 8'd16;
vramDataLower[12'd3921] = 8'd135;
vramDataLower[12'd3922] = 8'd90;
vramDataLower[12'd3923] = 8'd135;
vramDataLower[12'd3924] = 8'd166;
vramDataLower[12'd3925] = 8'd135;
vramDataLower[12'd3926] = 8'd202;
vramDataLower[12'd3927] = 8'd135;
vramDataLower[12'd3928] = 8'd31;
vramDataLower[12'd3929] = 8'd135;
vramDataLower[12'd3930] = 8'd202;
vramDataLower[12'd3931] = 8'd120;
vramDataLower[12'd3932] = 8'd16;
vramDataLower[12'd3933] = 8'd120;
vramDataLower[12'd3934] = 8'd202;
vramDataLower[12'd3935] = 8'd120;
vramDataLower[12'd3936] = 8'd202;
vramDataLower[12'd3937] = 8'd120;
vramDataLower[12'd3938] = 8'd75;
vramDataLower[12'd3939] = 8'd120;
vramDataLower[12'd3940] = 8'd31;
vramDataLower[12'd3941] = 8'd120;
vramDataLower[12'd3942] = 8'd16;
vramDataLower[12'd3943] = 8'd120;
vramDataLower[12'd3944] = 8'd145;
vramDataLower[12'd3945] = 8'd120;
vramDataLower[12'd3946] = 8'd52;
vramDataLower[12'd3947] = 8'd120;
vramDataLower[12'd3948] = 8'd30;
vramDataLower[12'd3949] = 8'd120;
vramDataLower[12'd3950] = 8'd17;
vramDataLower[12'd3951] = 8'd120;
vramDataLower[12'd3952] = 8'd198;
vramDataLower[12'd3953] = 8'd120;
vramDataLower[12'd3954] = 8'd145;
vramDataLower[12'd3955] = 8'd120;
vramDataLower[12'd3956] = 8'd164;
vramDataLower[12'd3957] = 8'd120;
vramDataLower[12'd3958] = 8'd83;
vramDataLower[12'd3959] = 8'd120;
vramDataLower[12'd3960] = 8'd83;
vramDataLower[12'd3961] = 8'd135;
vramDataLower[12'd3962] = 8'd30;
vramDataLower[12'd3963] = 8'd135;
vramDataLower[12'd3964] = 8'd37;
vramDataLower[12'd3965] = 8'd135;
vramDataLower[12'd3966] = 8'd62;
vramDataLower[12'd3967] = 8'd135;
vramDataLower[12'd3968] = 8'd61;
vramDataLower[12'd3969] = 8'd135;
vramDataLower[12'd3970] = 8'd94;
vramDataLower[12'd3971] = 8'd55;
vramDataLower[12'd3972] = 8'd46;
vramDataLower[12'd3973] = 8'd87;
vramDataLower[12'd3974] = 8'd214;
vramDataLower[12'd3975] = 8'd87;
vramDataLower[12'd3976] = 8'd28;
vramDataLower[12'd3977] = 8'd87;
vramDataLower[12'd3978] = 8'd0;
vramDataLower[12'd3979] = 8'd231;
vramDataLower[12'd3980] = 8'd252;
vramDataLower[12'd3981] = 8'd247;
vramDataLower[12'd3982] = 8'd183;
vramDataLower[12'd3983] = 8'd55;
vramDataLower[12'd3984] = 8'd255;
vramDataLower[12'd3985] = 8'd39;
vramDataLower[12'd3986] = 8'd198;
vramDataLower[12'd3987] = 8'd55;
vramDataLower[12'd3988] = 8'd202;
vramDataLower[12'd3989] = 8'd56;
vramDataLower[12'd3990] = 8'd223;
vramDataLower[12'd3991] = 8'd48;
vramDataLower[12'd3992] = 8'd223;
vramDataLower[12'd3993] = 8'd48;
vramDataLower[12'd3994] = 8'd223;
vramDataLower[12'd3995] = 8'd48;
vramDataLower[12'd3996] = 8'd223;
vramDataLower[12'd3997] = 8'd48;
vramDataLower[12'd3998] = 8'd220;
vramDataLower[12'd3999] = 8'd131;
vramDataLower[12'd4000] = 8'd210;
vramDataLower[12'd4001] = 8'd152;
vramDataLower[12'd4002] = 8'd164;
vramDataLower[12'd4003] = 8'd152;
vramDataLower[12'd4004] = 8'd210;
vramDataLower[12'd4005] = 8'd152;
vramDataLower[12'd4006] = 8'd210;
vramDataLower[12'd4007] = 8'd152;
vramDataLower[12'd4008] = 8'd145;
vramDataLower[12'd4009] = 8'd152;
vramDataLower[12'd4010] = 8'd145;
vramDataLower[12'd4011] = 8'd152;
vramDataLower[12'd4012] = 8'd48;
vramDataLower[12'd4013] = 8'd152;
vramDataLower[12'd4014] = 8'd148;
vramDataLower[12'd4015] = 8'd152;
vramDataLower[12'd4016] = 8'd202;
vramDataLower[12'd4017] = 8'd152;
vramDataLower[12'd4018] = 8'd164;
vramDataLower[12'd4019] = 8'd152;
vramDataLower[12'd4020] = 8'd210;
vramDataLower[12'd4021] = 8'd152;
vramDataLower[12'd4022] = 8'd181;
vramDataLower[12'd4023] = 8'd152;
vramDataLower[12'd4024] = 8'd198;
vramDataLower[12'd4025] = 8'd120;
vramDataLower[12'd4026] = 8'd210;
vramDataLower[12'd4027] = 8'd120;
vramDataLower[12'd4028] = 8'd16;
vramDataLower[12'd4029] = 8'd152;
vramDataLower[12'd4030] = 8'd202;
vramDataLower[12'd4031] = 8'd152;
vramDataLower[12'd4032] = 8'd164;
vramDataLower[12'd4033] = 8'd152;
vramDataLower[12'd4034] = 8'd50;
vramDataLower[12'd4035] = 8'd120;
vramDataLower[12'd4036] = 8'd190;
vramDataLower[12'd4037] = 8'd8;
vramDataLower[12'd4038] = 8'd139;
vramDataLower[12'd4039] = 8'd120;
vramDataLower[12'd4040] = 8'd92;
vramDataLower[12'd4041] = 8'd120;
vramDataLower[12'd4042] = 8'd198;
vramDataLower[12'd4043] = 8'd120;
vramDataLower[12'd4044] = 8'd135;
vramDataLower[12'd4045] = 8'd120;
vramDataLower[12'd4046] = 8'd200;
vramDataLower[12'd4047] = 8'd120;
vramDataLower[12'd4048] = 8'd172;
vramDataLower[12'd4049] = 8'd120;
vramDataLower[12'd4050] = 8'd31;
vramDataLower[12'd4051] = 8'd120;
vramDataLower[12'd4052] = 8'd16;
vramDataLower[12'd4053] = 8'd120;
vramDataLower[12'd4054] = 8'd183;
vramDataLower[12'd4055] = 8'd120;
vramDataLower[12'd4056] = 8'd183;
vramDataLower[12'd4057] = 8'd120;
vramDataLower[12'd4058] = 8'd164;
vramDataLower[12'd4059] = 8'd8;
vramDataLower[12'd4060] = 8'd16;
vramDataLower[12'd4061] = 8'd8;
vramDataLower[12'd4062] = 8'd70;
vramDataLower[12'd4063] = 8'd120;
vramDataLower[12'd4064] = 8'd200;
vramDataLower[12'd4065] = 8'd120;
vramDataLower[12'd4066] = 8'd155;
vramDataLower[12'd4067] = 8'd120;
vramDataLower[12'd4068] = 8'd202;
vramDataLower[12'd4069] = 8'd120;
vramDataLower[12'd4070] = 8'd228;
vramDataLower[12'd4071] = 8'd135;
vramDataLower[12'd4072] = 8'd210;
vramDataLower[12'd4073] = 8'd135;
vramDataLower[12'd4074] = 8'd37;
vramDataLower[12'd4075] = 8'd135;
vramDataLower[12'd4076] = 8'd183;
vramDataLower[12'd4077] = 8'd135;
vramDataLower[12'd4078] = 8'd202;
vramDataLower[12'd4079] = 8'd135;
vramDataLower[12'd4080] = 8'd230;
vramDataLower[12'd4081] = 8'd120;
vramDataLower[12'd4082] = 8'd16;
vramDataLower[12'd4083] = 8'd135;
vramDataLower[12'd4084] = 8'd50;
vramDataLower[12'd4085] = 8'd135;
vramDataLower[12'd4086] = 8'd135;
vramDataLower[12'd4087] = 8'd135;
vramDataLower[12'd4088] = 8'd85;
vramDataLower[12'd4089] = 8'd135;
vramDataLower[12'd4090] = 8'd17;
vramDataLower[12'd4091] = 8'd120;
vramDataLower[12'd4092] = 8'd156;
vramDataLower[12'd4093] = 8'd120;
vramDataLower[12'd4094] = 8'd90;
vramDataLower[12'd4095] = 8'd120;
