vramDataUpper[10'd0] = 8'd125;
vramDataUpper[10'd1] = 8'd120;
vramDataUpper[10'd2] = 8'd44;
vramDataUpper[10'd3] = 8'd120;
vramDataUpper[10'd4] = 8'd92;
vramDataUpper[10'd5] = 8'd120;
vramDataUpper[10'd6] = 8'd183;
vramDataUpper[10'd7] = 8'd120;
vramDataUpper[10'd8] = 8'd30;
vramDataUpper[10'd9] = 8'd120;
vramDataUpper[10'd10] = 8'd80;
vramDataUpper[10'd11] = 8'd120;
vramDataUpper[10'd12] = 8'd16;
vramDataUpper[10'd13] = 8'd120;
vramDataUpper[10'd14] = 8'd30;
vramDataUpper[10'd15] = 8'd120;
vramDataUpper[10'd16] = 8'd80;
vramDataUpper[10'd17] = 8'd135;
vramDataUpper[10'd18] = 8'd183;
vramDataUpper[10'd19] = 8'd120;
vramDataUpper[10'd20] = 8'd31;
vramDataUpper[10'd21] = 8'd120;
vramDataUpper[10'd22] = 8'd164;
vramDataUpper[10'd23] = 8'd120;
vramDataUpper[10'd24] = 8'd37;
vramDataUpper[10'd25] = 8'd120;
vramDataUpper[10'd26] = 8'd83;
vramDataUpper[10'd27] = 8'd135;
vramDataUpper[10'd28] = 8'd104;
vramDataUpper[10'd29] = 8'd135;
vramDataUpper[10'd30] = 8'd114;
vramDataUpper[10'd31] = 8'd135;
vramDataUpper[10'd32] = 8'd95;
vramDataUpper[10'd33] = 8'd135;
vramDataUpper[10'd34] = 8'd218;
vramDataUpper[10'd35] = 8'd135;
vramDataUpper[10'd36] = 8'd70;
vramDataUpper[10'd37] = 8'd135;
vramDataUpper[10'd38] = 8'd228;
vramDataUpper[10'd39] = 8'd135;
vramDataUpper[10'd40] = 8'd96;
vramDataUpper[10'd41] = 8'd87;
vramDataUpper[10'd42] = 8'd218;
vramDataUpper[10'd43] = 8'd55;
vramDataUpper[10'd44] = 8'd210;
vramDataUpper[10'd45] = 8'd135;
vramDataUpper[10'd46] = 8'd16;
vramDataUpper[10'd47] = 8'd135;
vramDataUpper[10'd48] = 8'd0;
vramDataUpper[10'd49] = 8'd167;
vramDataUpper[10'd50] = 8'd198;
vramDataUpper[10'd51] = 8'd135;
vramDataUpper[10'd52] = 8'd198;
vramDataUpper[10'd53] = 8'd8;
vramDataUpper[10'd54] = 8'd210;
vramDataUpper[10'd55] = 8'd128;
vramDataUpper[10'd56] = 8'd210;
vramDataUpper[10'd57] = 8'd16;
vramDataUpper[10'd58] = 8'd210;
vramDataUpper[10'd59] = 8'd16;
vramDataUpper[10'd60] = 8'd210;
vramDataUpper[10'd61] = 8'd16;
vramDataUpper[10'd62] = 8'd210;
vramDataUpper[10'd63] = 8'd16;
vramDataUpper[10'd64] = 8'd202;
vramDataUpper[10'd65] = 8'd152;
vramDataUpper[10'd66] = 8'd164;
vramDataUpper[10'd67] = 8'd152;
vramDataUpper[10'd68] = 8'd202;
vramDataUpper[10'd69] = 8'd152;
vramDataUpper[10'd70] = 8'd16;
vramDataUpper[10'd71] = 8'd152;
vramDataUpper[10'd72] = 8'd202;
vramDataUpper[10'd73] = 8'd152;
vramDataUpper[10'd74] = 8'd83;
vramDataUpper[10'd75] = 8'd152;
vramDataUpper[10'd76] = 8'd16;
vramDataUpper[10'd77] = 8'd152;
vramDataUpper[10'd78] = 8'd202;
vramDataUpper[10'd79] = 8'd152;
vramDataUpper[10'd80] = 8'd210;
vramDataUpper[10'd81] = 8'd152;
vramDataUpper[10'd82] = 8'd210;
vramDataUpper[10'd83] = 8'd120;
vramDataUpper[10'd84] = 8'd16;
vramDataUpper[10'd85] = 8'd120;
vramDataUpper[10'd86] = 8'd80;
vramDataUpper[10'd87] = 8'd120;
vramDataUpper[10'd88] = 8'd202;
vramDataUpper[10'd89] = 8'd120;
vramDataUpper[10'd90] = 8'd202;
vramDataUpper[10'd91] = 8'd120;
vramDataUpper[10'd92] = 8'd164;
vramDataUpper[10'd93] = 8'd152;
vramDataUpper[10'd94] = 8'd16;
vramDataUpper[10'd95] = 8'd152;
vramDataUpper[10'd96] = 8'd195;
vramDataUpper[10'd97] = 8'd8;
vramDataUpper[10'd98] = 8'd166;
vramDataUpper[10'd99] = 8'd152;
vramDataUpper[10'd100] = 8'd200;
vramDataUpper[10'd101] = 8'd120;
vramDataUpper[10'd102] = 8'd85;
vramDataUpper[10'd103] = 8'd120;
vramDataUpper[10'd104] = 8'd173;
vramDataUpper[10'd105] = 8'd120;
vramDataUpper[10'd106] = 8'd37;
vramDataUpper[10'd107] = 8'd120;
vramDataUpper[10'd108] = 8'd251;
vramDataUpper[10'd109] = 8'd120;
vramDataUpper[10'd110] = 8'd31;
vramDataUpper[10'd111] = 8'd120;
vramDataUpper[10'd112] = 8'd236;
vramDataUpper[10'd113] = 8'd120;
vramDataUpper[10'd114] = 8'd17;
vramDataUpper[10'd115] = 8'd120;
vramDataUpper[10'd116] = 8'd86;
vramDataUpper[10'd117] = 8'd8;
vramDataUpper[10'd118] = 8'd239;
vramDataUpper[10'd119] = 8'd8;
vramDataUpper[10'd120] = 8'd94;
vramDataUpper[10'd121] = 8'd120;
vramDataUpper[10'd122] = 8'd31;
vramDataUpper[10'd123] = 8'd120;
vramDataUpper[10'd124] = 8'd101;
vramDataUpper[10'd125] = 8'd120;
vramDataUpper[10'd126] = 8'd17;
vramDataUpper[10'd127] = 8'd120;
vramDataUpper[10'd128] = 8'd16;
vramDataUpper[10'd129] = 8'd120;
vramDataUpper[10'd130] = 8'd16;
vramDataUpper[10'd131] = 8'd120;
vramDataUpper[10'd132] = 8'd28;
vramDataUpper[10'd133] = 8'd120;
vramDataUpper[10'd134] = 8'd17;
vramDataUpper[10'd135] = 8'd120;
vramDataUpper[10'd136] = 8'd228;
vramDataUpper[10'd137] = 8'd120;
vramDataUpper[10'd138] = 8'd214;
vramDataUpper[10'd139] = 8'd120;
vramDataUpper[10'd140] = 8'd17;
vramDataUpper[10'd141] = 8'd135;
vramDataUpper[10'd142] = 8'd76;
vramDataUpper[10'd143] = 8'd135;
vramDataUpper[10'd144] = 8'd197;
vramDataUpper[10'd145] = 8'd135;
vramDataUpper[10'd146] = 8'd202;
vramDataUpper[10'd147] = 8'd120;
vramDataUpper[10'd148] = 8'd202;
vramDataUpper[10'd149] = 8'd120;
vramDataUpper[10'd150] = 8'd155;
vramDataUpper[10'd151] = 8'd120;
vramDataUpper[10'd152] = 8'd164;
vramDataUpper[10'd153] = 8'd120;
vramDataUpper[10'd154] = 8'd18;
vramDataUpper[10'd155] = 8'd120;
vramDataUpper[10'd156] = 8'd16;
vramDataUpper[10'd157] = 8'd120;
vramDataUpper[10'd158] = 8'd141;
vramDataUpper[10'd159] = 8'd120;
vramDataUpper[10'd160] = 8'd171;
vramDataUpper[10'd161] = 8'd120;
vramDataUpper[10'd162] = 8'd41;
vramDataUpper[10'd163] = 8'd120;
vramDataUpper[10'd164] = 8'd213;
vramDataUpper[10'd165] = 8'd120;
vramDataUpper[10'd166] = 8'd135;
vramDataUpper[10'd167] = 8'd120;
vramDataUpper[10'd168] = 8'd200;
vramDataUpper[10'd169] = 8'd120;
vramDataUpper[10'd170] = 8'd18;
vramDataUpper[10'd171] = 8'd120;
vramDataUpper[10'd172] = 8'd208;
vramDataUpper[10'd173] = 8'd120;
vramDataUpper[10'd174] = 8'd148;
vramDataUpper[10'd175] = 8'd120;
vramDataUpper[10'd176] = 8'd31;
vramDataUpper[10'd177] = 8'd120;
vramDataUpper[10'd178] = 8'd172;
vramDataUpper[10'd179] = 8'd135;
vramDataUpper[10'd180] = 8'd48;
vramDataUpper[10'd181] = 8'd135;
vramDataUpper[10'd182] = 8'd149;
vramDataUpper[10'd183] = 8'd120;
vramDataUpper[10'd184] = 8'd16;
vramDataUpper[10'd185] = 8'd135;
vramDataUpper[10'd186] = 8'd207;
vramDataUpper[10'd187] = 8'd135;
vramDataUpper[10'd188] = 8'd17;
vramDataUpper[10'd189] = 8'd135;
vramDataUpper[10'd190] = 8'd37;
vramDataUpper[10'd191] = 8'd135;
vramDataUpper[10'd192] = 8'd210;
vramDataUpper[10'd193] = 8'd135;
vramDataUpper[10'd194] = 8'd145;
vramDataUpper[10'd195] = 8'd135;
vramDataUpper[10'd196] = 8'd16;
vramDataUpper[10'd197] = 8'd135;
vramDataUpper[10'd198] = 8'd94;
vramDataUpper[10'd199] = 8'd135;
vramDataUpper[10'd200] = 8'd214;
vramDataUpper[10'd201] = 8'd135;
vramDataUpper[10'd202] = 8'd16;
vramDataUpper[10'd203] = 8'd135;
vramDataUpper[10'd204] = 8'd83;
vramDataUpper[10'd205] = 8'd135;
vramDataUpper[10'd206] = 8'd80;
vramDataUpper[10'd207] = 8'd135;
vramDataUpper[10'd208] = 8'd163;
vramDataUpper[10'd209] = 8'd119;
vramDataUpper[10'd210] = 8'd198;
vramDataUpper[10'd211] = 8'd135;
vramDataUpper[10'd212] = 8'd230;
vramDataUpper[10'd213] = 8'd152;
vramDataUpper[10'd214] = 8'd183;
vramDataUpper[10'd215] = 8'd152;
vramDataUpper[10'd216] = 8'd202;
vramDataUpper[10'd217] = 8'd8;
vramDataUpper[10'd218] = 8'd202;
vramDataUpper[10'd219] = 8'd8;
vramDataUpper[10'd220] = 8'd202;
vramDataUpper[10'd221] = 8'd8;
vramDataUpper[10'd222] = 8'd202;
vramDataUpper[10'd223] = 8'd8;
vramDataUpper[10'd224] = 8'd210;
vramDataUpper[10'd225] = 8'd152;
vramDataUpper[10'd226] = 8'd210;
vramDataUpper[10'd227] = 8'd152;
vramDataUpper[10'd228] = 8'd210;
vramDataUpper[10'd229] = 8'd152;
vramDataUpper[10'd230] = 8'd210;
vramDataUpper[10'd231] = 8'd152;
vramDataUpper[10'd232] = 8'd210;
vramDataUpper[10'd233] = 8'd152;
vramDataUpper[10'd234] = 8'd210;
vramDataUpper[10'd235] = 8'd152;
vramDataUpper[10'd236] = 8'd210;
vramDataUpper[10'd237] = 8'd152;
vramDataUpper[10'd238] = 8'd202;
vramDataUpper[10'd239] = 8'd152;
vramDataUpper[10'd240] = 8'd202;
vramDataUpper[10'd241] = 8'd152;
vramDataUpper[10'd242] = 8'd183;
vramDataUpper[10'd243] = 8'd8;
vramDataUpper[10'd244] = 8'd202;
vramDataUpper[10'd245] = 8'd152;
vramDataUpper[10'd246] = 8'd202;
vramDataUpper[10'd247] = 8'd152;
vramDataUpper[10'd248] = 8'd202;
vramDataUpper[10'd249] = 8'd152;
vramDataUpper[10'd250] = 8'd248;
vramDataUpper[10'd251] = 8'd152;
vramDataUpper[10'd252] = 8'd252;
vramDataUpper[10'd253] = 8'd152;
vramDataUpper[10'd254] = 8'd200;
vramDataUpper[10'd255] = 8'd152;
vramDataUpper[10'd256] = 8'd210;
vramDataUpper[10'd257] = 8'd152;
vramDataUpper[10'd258] = 8'd230;
vramDataUpper[10'd259] = 8'd152;
vramDataUpper[10'd260] = 8'd249;
vramDataUpper[10'd261] = 8'd8;
vramDataUpper[10'd262] = 8'd218;
vramDataUpper[10'd263] = 8'd8;
vramDataUpper[10'd264] = 8'd84;
vramDataUpper[10'd265] = 8'd152;
vramDataUpper[10'd266] = 8'd252;
vramDataUpper[10'd267] = 8'd152;
vramDataUpper[10'd268] = 8'd75;
vramDataUpper[10'd269] = 8'd120;
vramDataUpper[10'd270] = 8'd110;
vramDataUpper[10'd271] = 8'd152;
vramDataUpper[10'd272] = 8'd48;
vramDataUpper[10'd273] = 8'd152;
vramDataUpper[10'd274] = 8'd212;
vramDataUpper[10'd275] = 8'd8;
vramDataUpper[10'd276] = 8'd169;
vramDataUpper[10'd277] = 8'd8;
vramDataUpper[10'd278] = 8'd202;
vramDataUpper[10'd279] = 8'd152;
vramDataUpper[10'd280] = 8'd28;
vramDataUpper[10'd281] = 8'd120;
vramDataUpper[10'd282] = 8'd74;
vramDataUpper[10'd283] = 8'd120;
vramDataUpper[10'd284] = 8'd16;
vramDataUpper[10'd285] = 8'd120;
vramDataUpper[10'd286] = 8'd166;
vramDataUpper[10'd287] = 8'd8;
vramDataUpper[10'd288] = 8'd155;
vramDataUpper[10'd289] = 8'd8;
vramDataUpper[10'd290] = 8'd198;
vramDataUpper[10'd291] = 8'd152;
vramDataUpper[10'd292] = 8'd84;
vramDataUpper[10'd293] = 8'd120;
vramDataUpper[10'd294] = 8'd16;
vramDataUpper[10'd295] = 8'd135;
vramDataUpper[10'd296] = 8'd200;
vramDataUpper[10'd297] = 8'd135;
vramDataUpper[10'd298] = 8'd210;
vramDataUpper[10'd299] = 8'd135;
vramDataUpper[10'd300] = 8'd202;
vramDataUpper[10'd301] = 8'd120;
vramDataUpper[10'd302] = 8'd202;
vramDataUpper[10'd303] = 8'd120;
vramDataUpper[10'd304] = 8'd16;
vramDataUpper[10'd305] = 8'd120;
vramDataUpper[10'd306] = 8'd202;
vramDataUpper[10'd307] = 8'd120;
vramDataUpper[10'd308] = 8'd230;
vramDataUpper[10'd309] = 8'd120;
vramDataUpper[10'd310] = 8'd214;
vramDataUpper[10'd311] = 8'd120;
vramDataUpper[10'd312] = 8'd197;
vramDataUpper[10'd313] = 8'd120;
vramDataUpper[10'd314] = 8'd159;
vramDataUpper[10'd315] = 8'd120;
vramDataUpper[10'd316] = 8'd17;
vramDataUpper[10'd317] = 8'd120;
vramDataUpper[10'd318] = 8'd202;
vramDataUpper[10'd319] = 8'd152;
vramDataUpper[10'd320] = 8'd126;
vramDataUpper[10'd321] = 8'd120;
vramDataUpper[10'd322] = 8'd200;
vramDataUpper[10'd323] = 8'd120;
vramDataUpper[10'd324] = 8'd16;
vramDataUpper[10'd325] = 8'd120;
vramDataUpper[10'd326] = 8'd183;
vramDataUpper[10'd327] = 8'd120;
vramDataUpper[10'd328] = 8'd171;
vramDataUpper[10'd329] = 8'd120;
vramDataUpper[10'd330] = 8'd92;
vramDataUpper[10'd331] = 8'd120;
vramDataUpper[10'd332] = 8'd95;
vramDataUpper[10'd333] = 8'd120;
vramDataUpper[10'd334] = 8'd92;
vramDataUpper[10'd335] = 8'd120;
vramDataUpper[10'd336] = 8'd18;
vramDataUpper[10'd337] = 8'd120;
vramDataUpper[10'd338] = 8'd162;
vramDataUpper[10'd339] = 8'd120;
vramDataUpper[10'd340] = 8'd37;
vramDataUpper[10'd341] = 8'd135;
vramDataUpper[10'd342] = 8'd48;
vramDataUpper[10'd343] = 8'd135;
vramDataUpper[10'd344] = 8'd129;
vramDataUpper[10'd345] = 8'd135;
vramDataUpper[10'd346] = 8'd171;
vramDataUpper[10'd347] = 8'd135;
vramDataUpper[10'd348] = 8'd148;
vramDataUpper[10'd349] = 8'd135;
vramDataUpper[10'd350] = 8'd83;
vramDataUpper[10'd351] = 8'd135;
vramDataUpper[10'd352] = 8'd16;
vramDataUpper[10'd353] = 8'd135;
vramDataUpper[10'd354] = 8'd248;
vramDataUpper[10'd355] = 8'd135;
vramDataUpper[10'd356] = 8'd214;
vramDataUpper[10'd357] = 8'd135;
vramDataUpper[10'd358] = 8'd80;
vramDataUpper[10'd359] = 8'd120;
vramDataUpper[10'd360] = 8'd198;
vramDataUpper[10'd361] = 8'd120;
vramDataUpper[10'd362] = 8'd210;
vramDataUpper[10'd363] = 8'd120;
vramDataUpper[10'd364] = 8'd67;
vramDataUpper[10'd365] = 8'd135;
vramDataUpper[10'd366] = 8'd248;
vramDataUpper[10'd367] = 8'd135;
vramDataUpper[10'd368] = 8'd183;
vramDataUpper[10'd369] = 8'd119;
vramDataUpper[10'd370] = 8'd198;
vramDataUpper[10'd371] = 8'd135;
vramDataUpper[10'd372] = 8'd210;
vramDataUpper[10'd373] = 8'd152;
vramDataUpper[10'd374] = 8'd210;
vramDataUpper[10'd375] = 8'd152;
vramDataUpper[10'd376] = 8'd210;
vramDataUpper[10'd377] = 8'd152;
vramDataUpper[10'd378] = 8'd210;
vramDataUpper[10'd379] = 8'd152;
vramDataUpper[10'd380] = 8'd210;
vramDataUpper[10'd381] = 8'd24;
vramDataUpper[10'd382] = 8'd31;
vramDataUpper[10'd383] = 8'd152;
vramDataUpper[10'd384] = 8'd210;
vramDataUpper[10'd385] = 8'd152;
vramDataUpper[10'd386] = 8'd164;
vramDataUpper[10'd387] = 8'd152;
vramDataUpper[10'd388] = 8'd209;
vramDataUpper[10'd389] = 8'd152;
vramDataUpper[10'd390] = 8'd164;
vramDataUpper[10'd391] = 8'd152;
vramDataUpper[10'd392] = 8'd83;
vramDataUpper[10'd393] = 8'd152;
vramDataUpper[10'd394] = 8'd181;
vramDataUpper[10'd395] = 8'd152;
vramDataUpper[10'd396] = 8'd80;
vramDataUpper[10'd397] = 8'd152;
vramDataUpper[10'd398] = 8'd210;
vramDataUpper[10'd399] = 8'd8;
vramDataUpper[10'd400] = 8'd210;
vramDataUpper[10'd401] = 8'd8;
vramDataUpper[10'd402] = 8'd183;
vramDataUpper[10'd403] = 8'd8;
vramDataUpper[10'd404] = 8'd90;
vramDataUpper[10'd405] = 8'd8;
vramDataUpper[10'd406] = 8'd17;
vramDataUpper[10'd407] = 8'd152;
vramDataUpper[10'd408] = 8'd248;
vramDataUpper[10'd409] = 8'd152;
vramDataUpper[10'd410] = 8'd209;
vramDataUpper[10'd411] = 8'd8;
vramDataUpper[10'd412] = 8'd210;
vramDataUpper[10'd413] = 8'd8;
vramDataUpper[10'd414] = 8'd183;
vramDataUpper[10'd415] = 8'd8;
vramDataUpper[10'd416] = 8'd212;
vramDataUpper[10'd417] = 8'd152;
vramDataUpper[10'd418] = 8'd31;
vramDataUpper[10'd419] = 8'd152;
vramDataUpper[10'd420] = 8'd210;
vramDataUpper[10'd421] = 8'd152;
vramDataUpper[10'd422] = 8'd210;
vramDataUpper[10'd423] = 8'd152;
vramDataUpper[10'd424] = 8'd135;
vramDataUpper[10'd425] = 8'd152;
vramDataUpper[10'd426] = 8'd166;
vramDataUpper[10'd427] = 8'd8;
vramDataUpper[10'd428] = 8'd95;
vramDataUpper[10'd429] = 8'd120;
vramDataUpper[10'd430] = 8'd250;
vramDataUpper[10'd431] = 8'd8;
vramDataUpper[10'd432] = 8'd124;
vramDataUpper[10'd433] = 8'd152;
vramDataUpper[10'd434] = 8'd95;
vramDataUpper[10'd435] = 8'd152;
vramDataUpper[10'd436] = 8'd210;
vramDataUpper[10'd437] = 8'd152;
vramDataUpper[10'd438] = 8'd106;
vramDataUpper[10'd439] = 8'd120;
vramDataUpper[10'd440] = 8'd214;
vramDataUpper[10'd441] = 8'd120;
vramDataUpper[10'd442] = 8'd210;
vramDataUpper[10'd443] = 8'd120;
vramDataUpper[10'd444] = 8'd210;
vramDataUpper[10'd445] = 8'd120;
vramDataUpper[10'd446] = 8'd202;
vramDataUpper[10'd447] = 8'd135;
vramDataUpper[10'd448] = 8'd16;
vramDataUpper[10'd449] = 8'd135;
vramDataUpper[10'd450] = 8'd109;
vramDataUpper[10'd451] = 8'd120;
vramDataUpper[10'd452] = 8'd31;
vramDataUpper[10'd453] = 8'd120;
vramDataUpper[10'd454] = 8'd171;
vramDataUpper[10'd455] = 8'd120;
vramDataUpper[10'd456] = 8'd83;
vramDataUpper[10'd457] = 8'd120;
vramDataUpper[10'd458] = 8'd230;
vramDataUpper[10'd459] = 8'd120;
vramDataUpper[10'd460] = 8'd90;
vramDataUpper[10'd461] = 8'd120;
vramDataUpper[10'd462] = 8'd16;
vramDataUpper[10'd463] = 8'd120;
vramDataUpper[10'd464] = 8'd159;
vramDataUpper[10'd465] = 8'd120;
vramDataUpper[10'd466] = 8'd17;
vramDataUpper[10'd467] = 8'd120;
vramDataUpper[10'd468] = 8'd202;
vramDataUpper[10'd469] = 8'd120;
vramDataUpper[10'd470] = 8'd16;
vramDataUpper[10'd471] = 8'd120;
vramDataUpper[10'd472] = 8'd166;
vramDataUpper[10'd473] = 8'd120;
vramDataUpper[10'd474] = 8'd16;
vramDataUpper[10'd475] = 8'd152;
vramDataUpper[10'd476] = 8'd28;
vramDataUpper[10'd477] = 8'd152;
vramDataUpper[10'd478] = 8'd28;
vramDataUpper[10'd479] = 8'd8;
vramDataUpper[10'd480] = 8'd209;
vramDataUpper[10'd481] = 8'd136;
vramDataUpper[10'd482] = 8'd39;
vramDataUpper[10'd483] = 8'd152;
vramDataUpper[10'd484] = 8'd80;
vramDataUpper[10'd485] = 8'd152;
vramDataUpper[10'd486] = 8'd200;
vramDataUpper[10'd487] = 8'd120;
vramDataUpper[10'd488] = 8'd31;
vramDataUpper[10'd489] = 8'd120;
vramDataUpper[10'd490] = 8'd17;
vramDataUpper[10'd491] = 8'd120;
vramDataUpper[10'd492] = 8'd30;
vramDataUpper[10'd493] = 8'd120;
vramDataUpper[10'd494] = 8'd17;
vramDataUpper[10'd495] = 8'd120;
vramDataUpper[10'd496] = 8'd135;
vramDataUpper[10'd497] = 8'd135;
vramDataUpper[10'd498] = 8'd90;
vramDataUpper[10'd499] = 8'd135;
vramDataUpper[10'd500] = 8'd83;
vramDataUpper[10'd501] = 8'd135;
vramDataUpper[10'd502] = 8'd30;
vramDataUpper[10'd503] = 8'd135;
vramDataUpper[10'd504] = 8'd202;
vramDataUpper[10'd505] = 8'd120;
vramDataUpper[10'd506] = 8'd210;
vramDataUpper[10'd507] = 8'd120;
vramDataUpper[10'd508] = 8'd80;
vramDataUpper[10'd509] = 8'd135;
vramDataUpper[10'd510] = 8'd172;
vramDataUpper[10'd511] = 8'd135;
vramDataUpper[10'd512] = 8'd210;
vramDataUpper[10'd513] = 8'd135;
vramDataUpper[10'd514] = 8'd80;
vramDataUpper[10'd515] = 8'd120;
vramDataUpper[10'd516] = 8'd75;
vramDataUpper[10'd517] = 8'd120;
vramDataUpper[10'd518] = 8'd202;
vramDataUpper[10'd519] = 8'd120;
vramDataUpper[10'd520] = 8'd90;
vramDataUpper[10'd521] = 8'd120;
vramDataUpper[10'd522] = 8'd135;
vramDataUpper[10'd523] = 8'd135;
vramDataUpper[10'd524] = 8'd202;
vramDataUpper[10'd525] = 8'd135;
vramDataUpper[10'd526] = 8'd76;
vramDataUpper[10'd527] = 8'd135;
vramDataUpper[10'd528] = 8'd183;
vramDataUpper[10'd529] = 8'd55;
vramDataUpper[10'd530] = 8'd198;
vramDataUpper[10'd531] = 8'd135;
vramDataUpper[10'd532] = 8'd145;
vramDataUpper[10'd533] = 8'd152;
vramDataUpper[10'd534] = 8'd210;
vramDataUpper[10'd535] = 8'd152;
vramDataUpper[10'd536] = 8'd210;
vramDataUpper[10'd537] = 8'd152;
vramDataUpper[10'd538] = 8'd202;
vramDataUpper[10'd539] = 8'd152;
vramDataUpper[10'd540] = 8'd210;
vramDataUpper[10'd541] = 8'd152;
vramDataUpper[10'd542] = 8'd16;
vramDataUpper[10'd543] = 8'd152;
vramDataUpper[10'd544] = 8'd202;
vramDataUpper[10'd545] = 8'd152;
vramDataUpper[10'd546] = 8'd210;
vramDataUpper[10'd547] = 8'd152;
vramDataUpper[10'd548] = 8'd210;
vramDataUpper[10'd549] = 8'd152;
vramDataUpper[10'd550] = 8'd16;
vramDataUpper[10'd551] = 8'd152;
vramDataUpper[10'd552] = 8'd202;
vramDataUpper[10'd553] = 8'd152;
vramDataUpper[10'd554] = 8'd202;
vramDataUpper[10'd555] = 8'd152;
vramDataUpper[10'd556] = 8'd30;
vramDataUpper[10'd557] = 8'd24;
vramDataUpper[10'd558] = 8'd202;
vramDataUpper[10'd559] = 8'd8;
vramDataUpper[10'd560] = 8'd80;
vramDataUpper[10'd561] = 8'd8;
vramDataUpper[10'd562] = 8'd80;
vramDataUpper[10'd563] = 8'd8;
vramDataUpper[10'd564] = 8'd183;
vramDataUpper[10'd565] = 8'd24;
vramDataUpper[10'd566] = 8'd214;
vramDataUpper[10'd567] = 8'd8;
vramDataUpper[10'd568] = 8'd210;
vramDataUpper[10'd569] = 8'd8;
vramDataUpper[10'd570] = 8'd210;
vramDataUpper[10'd571] = 8'd8;
vramDataUpper[10'd572] = 8'd202;
vramDataUpper[10'd573] = 8'd8;
vramDataUpper[10'd574] = 8'd210;
vramDataUpper[10'd575] = 8'd8;
vramDataUpper[10'd576] = 8'd83;
vramDataUpper[10'd577] = 8'd8;
vramDataUpper[10'd578] = 8'd183;
vramDataUpper[10'd579] = 8'd8;
vramDataUpper[10'd580] = 8'd210;
vramDataUpper[10'd581] = 8'd8;
vramDataUpper[10'd582] = 8'd230;
vramDataUpper[10'd583] = 8'd8;
vramDataUpper[10'd584] = 8'd207;
vramDataUpper[10'd585] = 8'd120;
vramDataUpper[10'd586] = 8'd16;
vramDataUpper[10'd587] = 8'd120;
vramDataUpper[10'd588] = 8'd85;
vramDataUpper[10'd589] = 8'd120;
vramDataUpper[10'd590] = 8'd230;
vramDataUpper[10'd591] = 8'd120;
vramDataUpper[10'd592] = 8'd16;
vramDataUpper[10'd593] = 8'd120;
vramDataUpper[10'd594] = 8'd80;
vramDataUpper[10'd595] = 8'd120;
vramDataUpper[10'd596] = 8'd80;
vramDataUpper[10'd597] = 8'd120;
vramDataUpper[10'd598] = 8'd202;
vramDataUpper[10'd599] = 8'd120;
vramDataUpper[10'd600] = 8'd31;
vramDataUpper[10'd601] = 8'd120;
vramDataUpper[10'd602] = 8'd202;
vramDataUpper[10'd603] = 8'd120;
vramDataUpper[10'd604] = 8'd80;
vramDataUpper[10'd605] = 8'd120;
vramDataUpper[10'd606] = 8'd70;
vramDataUpper[10'd607] = 8'd120;
vramDataUpper[10'd608] = 8'd202;
vramDataUpper[10'd609] = 8'd120;
vramDataUpper[10'd610] = 8'd80;
vramDataUpper[10'd611] = 8'd120;
vramDataUpper[10'd612] = 8'd208;
vramDataUpper[10'd613] = 8'd120;
vramDataUpper[10'd614] = 8'd183;
vramDataUpper[10'd615] = 8'd8;
vramDataUpper[10'd616] = 8'd83;
vramDataUpper[10'd617] = 8'd120;
vramDataUpper[10'd618] = 8'd179;
vramDataUpper[10'd619] = 8'd8;
vramDataUpper[10'd620] = 8'd95;
vramDataUpper[10'd621] = 8'd8;
vramDataUpper[10'd622] = 8'd34;
vramDataUpper[10'd623] = 8'd120;
vramDataUpper[10'd624] = 8'd252;
vramDataUpper[10'd625] = 8'd120;
vramDataUpper[10'd626] = 8'd16;
vramDataUpper[10'd627] = 8'd120;
vramDataUpper[10'd628] = 8'd252;
vramDataUpper[10'd629] = 8'd152;
vramDataUpper[10'd630] = 8'd94;
vramDataUpper[10'd631] = 8'd152;
vramDataUpper[10'd632] = 8'd191;
vramDataUpper[10'd633] = 8'd152;
vramDataUpper[10'd634] = 8'd166;
vramDataUpper[10'd635] = 8'd152;
vramDataUpper[10'd636] = 8'd34;
vramDataUpper[10'd637] = 8'd152;
vramDataUpper[10'd638] = 8'd94;
vramDataUpper[10'd639] = 8'd152;
vramDataUpper[10'd640] = 8'd248;
vramDataUpper[10'd641] = 8'd152;
vramDataUpper[10'd642] = 8'd17;
vramDataUpper[10'd643] = 8'd120;
vramDataUpper[10'd644] = 8'd31;
vramDataUpper[10'd645] = 8'd152;
vramDataUpper[10'd646] = 8'd7;
vramDataUpper[10'd647] = 8'd120;
vramDataUpper[10'd648] = 8'd16;
vramDataUpper[10'd649] = 8'd152;
vramDataUpper[10'd650] = 8'd95;
vramDataUpper[10'd651] = 8'd120;
vramDataUpper[10'd652] = 8'd202;
vramDataUpper[10'd653] = 8'd120;
vramDataUpper[10'd654] = 8'd30;
vramDataUpper[10'd655] = 8'd120;
vramDataUpper[10'd656] = 8'd17;
vramDataUpper[10'd657] = 8'd120;
vramDataUpper[10'd658] = 8'd198;
vramDataUpper[10'd659] = 8'd120;
vramDataUpper[10'd660] = 8'd135;
vramDataUpper[10'd661] = 8'd120;
vramDataUpper[10'd662] = 8'd16;
vramDataUpper[10'd663] = 8'd135;
vramDataUpper[10'd664] = 8'd210;
vramDataUpper[10'd665] = 8'd135;
vramDataUpper[10'd666] = 8'd80;
vramDataUpper[10'd667] = 8'd120;
vramDataUpper[10'd668] = 8'd188;
vramDataUpper[10'd669] = 8'd120;
vramDataUpper[10'd670] = 8'd252;
vramDataUpper[10'd671] = 8'd120;
vramDataUpper[10'd672] = 8'd76;
vramDataUpper[10'd673] = 8'd152;
vramDataUpper[10'd674] = 8'd31;
vramDataUpper[10'd675] = 8'd120;
vramDataUpper[10'd676] = 8'd164;
vramDataUpper[10'd677] = 8'd152;
vramDataUpper[10'd678] = 8'd30;
vramDataUpper[10'd679] = 8'd120;
vramDataUpper[10'd680] = 8'd202;
vramDataUpper[10'd681] = 8'd120;
vramDataUpper[10'd682] = 8'd80;
vramDataUpper[10'd683] = 8'd120;
vramDataUpper[10'd684] = 8'd252;
vramDataUpper[10'd685] = 8'd120;
vramDataUpper[10'd686] = 8'd16;
vramDataUpper[10'd687] = 8'd135;
vramDataUpper[10'd688] = 8'd210;
vramDataUpper[10'd689] = 8'd135;
vramDataUpper[10'd690] = 8'd51;
vramDataUpper[10'd691] = 8'd135;
vramDataUpper[10'd692] = 8'd164;
vramDataUpper[10'd693] = 8'd152;
vramDataUpper[10'd694] = 8'd202;
vramDataUpper[10'd695] = 8'd152;
vramDataUpper[10'd696] = 8'd210;
vramDataUpper[10'd697] = 8'd152;
vramDataUpper[10'd698] = 8'd210;
vramDataUpper[10'd699] = 8'd152;
vramDataUpper[10'd700] = 8'd164;
vramDataUpper[10'd701] = 8'd152;
vramDataUpper[10'd702] = 8'd210;
vramDataUpper[10'd703] = 8'd152;
